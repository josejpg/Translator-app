Vanliga kommandoknappar  
Avbryt  
När du avslutar en dialogruta med kommandoknappen Avbryt stängs dialogen utan att de gjorda ändringarna övertas.  
Utrullningslist  
En del ikoner öppnar utrullningslister när man klickar på dem.  
Det är menyer där du kan välja bland olika element genom att klicka med musen.  
Men du kan också flytta hela utrullningslisten med musen om du pekar på titellisten, trycker på musknappen och håller ner den samtidigt som du drar den bort från sin plats.  
När du släpper musknappen stannar utrullningslisten på det nya stället.  
Du kan sedan flytta den genom att ta tag i titellisten och dra den till ett annat ställe eller stänga den genom att klicka på stäng-fönstret-symbolen.  
Rotationsfält  
Ange det numeriska värdet i det här textfältet eller välj det med pil-uppåt - eller pil-nedåt-knapparna.  
Du ställer in det maximala och minimala värdet för rotationsfältet med Page Up och Page Down.  
Om det rör sig om ett rotationsfält för numeriska värden kan du också ange en måttenhet, t.ex. 1 cm eller 5 mm eller 12 pt eller 2" (för 2 tum).  
Konvertera  
Om du klickar dig framåt genom dialogrutan, heter den här kommandoknappen Nästa>>.  
På sista sidan ändrar den namn till Konvertera.  
Om du klickar på kommandoknappen genomförs konverteringen.  
Snabbmeny  
Håll sedan ner Ctrl-tangenten respektive kommando - och alternativtangenten och klicka med musknappen höger musknapp på objektet. (Till en del objekt kan du också öppna snabbmenyn utan att först markera objektet.) Snabbmenyer finns nästan överallt i %PRODUCTNAME.  
Radera...  
Raderar det eller de markerade elementen efter en kontrollfråga.  
Radera  
Raderar det eller de markerade elementen utan någon kontrollfråga.  
Metrik  
I inmatningsfälten kan du ange värden i olika måttenheter.  
Standardmåttenheten är centimeter.  
Om du vill att avståndet t.ex. ska vara exakt 1 tum skriver du "1".  
Beroende på sammanhanget är fler enheter möjliga, t.ex. 12 pt för ett avstånd på 12 punkter.  
Om värdet är orealistiskt byter programmet ut det mot ett eget maximi - eller minimivärde.  
Stäng  
Med denna kommandoknapp stänger Du dialogrutan och alla ändringar som gjorts i dialogrutan övertas.  
Stäng  
Med denna kommandoknapp stänger Du dialogrutan.  
Standard  
Återställer de värden som visas i dialogrutan till de förinmatade standardvärdena, i den mån Du som användare kan påverka värdena.  
Det Du matar in som alternativ där har företräde framför programmets "fabriksinställningar", som gäller under installationen.  
Du får ingen kontrollfråga innan värdena återställs till standardvärdena.  
Om Du därefter bekräftar dialogrutan har de ändringar som Du gjort oåterkalleligen gått förlorade.  
Överta  
Övertar ändrade eller markerade värden utan att stänga dialogrutan.  
Förminska / förstora  
Klicka på den här symbolen om Du vill förminska dialogrutan så att den blir lika stor som inmatningsfältet eller för att återställa den till den ursprungliga storleken.  
Det blir då enklare att markera den önskade referensen i tabellen.  
Symbolen blir automatiskt en förstora-symbol.  
Klicka på ikonen Förstora, varpå dialogrutan återställs.  
Dialogrutan förminskas automatiskt om Du klickar med musknappen i tabellen och skapar ett område.  
Så snart Du släpper upp musknappen återgår dialogrutan till full storlek och den områdesreferens som definierats med musen markeras med en blå ram i dokumentet.  
Förminska  
Förstora  
Förhandsvisningsfält  
I detta fält ser Du hur de ändringar som Du nu kan utföra kommer att påverka dokumentet.  
Ett stiliserat exempel visas.  
Nästa  
När Du klickar på den här knappen använder AutoPiloten de aktuella inställningarna i dialogrutan och går vidare till nästa redigeringssteg.  
När Du kommit till det sista steget kallas denna kommandoknapp för Färdigställ.  
Tillbaka  
Återställer ändrade värden till standardvärdena.  
Det är de värden som gällde när applikationen öppnades.  
Du får ingen kontrollfråga innan värdena återställs till standardvärdena.  
Om Du därefter bekräftar dialogrutan har de ändringar som Du gjort oåterkalleligen gått förlorade.  
Tillbaka  
Återställer de ändringar som gjorts under den aktuella fliken till de inställningar som gällde när fliken öppnades.  
Någon kontrollfråga visas inte.  
Tillbaka  
I dialogrutan kan Du visa Dina val från det föregående arbetssteget.  
Aktuella inställningar bibehålls.  
Denna kommandoknapp är endast tillgänglig fr o m andra redigeringssteget.  
Återställ  
Återställer ändrade värden till standardvärdena.  
Du får ingen kontrollfråga innan värdena återställs till standardvärdena.  
Om Du därefter bekräftar dialogrutan har de ändringar som Du gjort oåterkalleligen gått förlorade.  
Fler  
Genom att klicka på denna kommandoknapp utvidgar Du dialogrutan med ytterligare alternativ.  
Genom att klicka en gång till återställer Du dialogrutans ursprungliga vy.  
Se även följande funktioner:  
Den här funktionen finns bara med om du har installerat analysadd-in.  
Sökningen stöder reguljära uttryck.  
Så snart du skriver in en söktext kan du t.ex. ange all* om du vill komma till den första sökträffen där tecknen "all" står åtföljda av godtyckliga tecken.  
Vid fel returnerar funktionen ett logiskt eller ett numeriskt värde.  
(Det här kommandot är bara tillgängligt via snabbmenyn).  
Du kan dubbelklicka på alla verktyg om du vill välja det som nytt verktyg permanent.  
Då kan du kan t.ex. rita ett flertal rektanglar efter varandra, tills du väljer ett nytt verktyg.  
Men om du bara aktiverar ett verktyg genom att klicka en gång på det, används det bara en gång, d.v.s. tills du t.ex. ritat klart den första rektangeln.  
Därefter växlar programmet automatiskt tillbaka till det tidigare valda verktyget.  
Facktermer enkelt förklarade - Internet-ordlista  
För att det ska bli lättare för dig att komma igång, finns här en ordlista som innehåller förklaringar av de viktigaste facktermerna inom områdena Internet, intranät, e-post och nyheter.  
Om du är nykomling på Internet stöter du säkert på många nya ord, som t.ex. browser, bookmark, e-mail, hemsida, sökmotor.  
Här får du reda på vad de här termerna och många andra betyder.  
Klicka på termen eller bläddra igenom förklaringen.  
applet, bookmark, browser, e-mail, frame (ram), FTP, HTML, HTTP, hyperlink, image map, intranet, Java, plug-in, proxy, server, SGML, SMTP / POP3, style sheet, sökmotor, tag, TCP / IP, URL, Web server, XML  
Applet  
Med applet (appletprogram) menar man på Internet-språk ett speciellt objekt som finns på en HTML -sida.  
Det innehåller ett program som är skrivet på Java, det mest använda språket på Internet.  
Animationen laddas inte som en rad enskilda bilder (som på en filmrulle) via Internet utan som ett program som körs i din webbläsare.  
Appletprogram kan användas till animationer, animerade texter, interaktiv inmatning av användaruppgifter, spel mm.  
I %PRODUCTNAME kan du infoga appletprogram som du själv har utvecklat eller laddat ner från Internet på dina sidor (menykommandot Infoga - Objekt - Applet).  
Sådana objekt kan sedan ses av alla användare som har en webbläsare som kan köra dina appletprogram.  
Webbläsare som inte klarar av det hoppar som regel bara över appletprogrammen.  
Du hittar många exempel på appletprogram på adressen http: / /www.gamelan.com.  
Bookmark  
I %PRODUCTNAME kan du sätta ett bokmärke till den aktuella hjälpsidan i hjälpfönstret.  
Browser  
Det kan användas t.ex. vid sökning av viss information.  
E-mail  
E-mail står för Electronic Mail (elektronisk post; e-post) och är meddelanden som skickas i ett kommunikationssystem, som t.ex. Internet.  
E-post kan innehålla information i form av text, bilder, ljud och andra bifogade filer.  
I %PRODUCTNAME kan du t.ex. skicka det aktuella dokumentet under Arkiv - Skicka som bilaga till ett e-brev.  
Då öppnas ditt standardprogram för e-post.  
Frame (ram)  
Frames (ramar) är en viktig del i layouten av HTML -sidor.  
I %PRODUCTNAME kan du använda fria ramar (floating frames).  
Ramar kan innehålla objekt, t.ex. grafik, videofiler och ljud, och kan infogas på HMTL-sidor.  
Några av dessa alternativ finns även på menyn Redigera - Objekt när ramen är markerad.  
FTP  
FTP står för File Transfer Protocol (protokoll för filöverföring) och är det normala överföringsprotokollet för filer på Internet.  
På den här datorn lagras filer som kan överföras med FTP.  
Medan FTP alltså är avsett för överföring och "nedladdning" av filer på Internet, är protokollet HTTP (Hypertext Transfer Protocol) till för uppkoppling och datautbyte mellan WWW-servrar och WWW-klienter.  
HTML  
HTML (Hypertext Markup Language) är ett dokumentbeskrivningsspråk som används som filformat för WWW-dokument.  
Det har sitt ursprung i SGML och kan hantera text, grafik, video och ljud.  
HTML (utförlig förklaring).  
HTML (utförlig förklaring)  
Om du vill skriva in HTML-kommandon direkt (t.ex. när du gör övningsuppgifterna i någon av de många HTML-handböcker som finns), måste du tänka på att HTML-sidor är rena textfiler i 7-bitars ASCII -kod.  
Spara alltså de dokument som du skriver direkt i HTML-kod och utan omljud (t.ex. å, ä, ö) och andra specialtecken i den utökade teckenuppsättningen som dokumenttypen Text DOS.  
Ge dem filnamnstillägget .HTM.  
Om du vill öppna den här filen i %PRODUCTNAME senare och fortsätta att redigera HTML-koden, måste du ladda den med filtypen Text DOS, inte med filtypen Webbsida.  
Det finns en mycket bra introduktion till HTML på svenska på http: / /www.skolverket.se / skolnet / htmlkurs /.  
HTTP  
Överföringsprotokollet för hypertext (HyperText Transfer Protocol) används för WWW-dokument mellan WWW - servrar (hosts) och webbläsare (klienter).  
Hyperlink  
Du kan aktivera dessa hänvisningar genom att klicka på dem.  
Med hjälp av hyperlänkar kan läsaren av ett dokument hoppa till relaterad information i samma dokument eller i andra dokument.  
På Internet är det t.ex. vanligt att skapa hyperlänkar på den egna hemsidan som leder till andra webbplatser.  
I %PRODUCTNAME kan hyperlänkar tilldelas såväl text (se hyperlänklisten) som grafik och textramar (se fliken Hyperlänk i dialogrutan för grafik / ram / objekt och menyn Redigera - Image map).  
Image map  
En image map är ett grafikobjekt eller en textram med en länk.  
Du kan klicka på specifika områden på grafikobjektet respektive textramen, och kommer då till det mål, eller den URL, som området är länkat med.  
Själva områdena, liksom de länkade webbadresserna och texterna som ska visas när muspekaren pekar på något av områdena, definierar du i Image map-redigeraren.  
Det finns två image map-typer.  
Den ena typen, Client Side ImageMap, utvärderas av den måldator som har laddat grafikobjektet via Internet, medan den andra typen, Server Side ImageMap, utvärderas av den dator som tillhandahåller HTML -sidan på Internet.  
Vid serverutvärdering skickas markörens position på bilden eller ramen i relativa koordinater till servern när användaren klickar på en image map och ett särskilt program på servern reagerar utifrån denna information.  
Om du använder "modern" klientutvärdering och klickar på en definierad "hot spot "på en image map hämtas den därtill knutna URL-adressen, precis som om du hade klickat på en vanlig textlänk.  
Dessutom visas URL-adressen nedanför muspekaren när du pekar på bilden.  
Den här annorlunda funktionaliteten visar att image maps kan förekomma i mycket olika format.  
Image map-format  
De olika image map -typerna skiljer sig framför allt åt i ett avseende, nämligen om de utvärderas på servern (t.ex. hos Internet-leverantören) eller i webbläsaren på din egen dator.  
Image map på serversidan  
Image maps på servern visas som bilder eller ramar hos läsaren där han / hon kan klicka på dem med musen.  
Koordinaterna för muspekarens relativa position skickas till servern där ett särskilt program tar reda på vilken nästa åtgärd ska vara.  
Det finns flera metoder för att definiera detta förfaringssätt och de är inte kompatibla sinsemellan.  
De två vanligaste är:  
W3C (CERN) HTTP-server (formattyp:  
MAP - CERN)  
NCSA HTTP-server (formattyp:  
MAP - NCSA)  
Med %PRODUCTNAME kan du skapa image maps för båda metoderna.  
Du väljer format i listrutan Filtyp i dialogrutan Spara image map som.  
Separata map-filer skapas som du måste skicka till servern.  
Under alla omständigheter måste du fråga din Internetleverantör eller nätadministratör vilken typ av image map som stöds av servern och hur utvärderingsprogrammet ska "tilltalas".  
Image map på klientsidan  
Moderna image maps på klientdatorn kräver inte så stor insats av servern.  
Det område som läsaren kan klicka på i en bild eller en ram indikeras direkt när du pekar på det genom att den länkade URL -adressen visas.  
En image map ligger så att säga i ett skikt ovanför bilden och innehåller information om de klickbara områdena.  
Detta är dock något som får mindre betydelse allteftersom de äldre webbläsarna ersätts med nyare versioner.  
Om du väljer filtypen SIP - Starview ImageMap när du sparar en image map, lagras den automatiskt i ett format som gör att du kan använda den för alla grafikobjekt eller ramar som du har aktiverat i dokumentet.  
Däremot ska du inte spara en image map separat om du bara vill använda den för det aktuella grafikobjektet eller textramen.  
När du har definierat områdena klickar du på ikonen Tilldela.  
Mer behöver du inte göra.  
Image maps på klientdatorn infogas direkt i sidans HTML-kod när du sparar dem i HTML -format.  
Vissa mycket använda webbläsare utvärderar image maps på klientdatorn bildpunkt per bildpunkt så som de beskrivs i dokumentet.  
I %PRODUCTNAME beräknas storlekarna utifrån grafikobjektets originalstorlek och skalas vid träfftestet.  
För grafik med fasta storleksuppgifter och helt utan storleksuppgifter omräknas detta.  
För grafik med relativa storleksuppgifter används originalstorleken.  
Grafik med procentuella uppgifter behandlas av vissa andra webbläsare på ett felaktigt sätt, medan %PRODUCTNAME enbart visar användbara resultat.  
Intranät  
Ett intranät är ett lokalt nätverk som används för TCP / IP -kommunikation med överföringsprotokollet HTTP.  
Gentemot vanliga nätverk har ett intranät fördelen att det är mycket enkelt att övergå till Internet och att programvaran är mycket prisvärd för närvarande.  
IP-adress  
Den skrivs ut som fyra heltal mellan 0 och 255.  
Exempel:  
Varje användare har en sådan Internet-protokolladress.  
Ofta blir IP-adressen bara dynamiskt tilldelad och gäller alltså bara för den aktuella uppkopplingen.  
Eftersom det är krångligt att komma ihåg eller skriva ner den här typen av adresser, adresseras nästan alltid servrar på Internet enbart med sina namn.  
En dator som kallas namnserver ser till att namnet byts ut mot korrekt IP-adress.  
Java  
Java är ett s.k. plattformsoberoende (d.v.s. oberoende av operativsystem, processor mm) programmeringsspråk, utvecklat av Sun Microsystems, Inc (http: / /www.sun.com och http: / /www.sun.se).  
Webbsidor och tillämpningar som är programmerade med Java kan användas av alla plattformar som stöder detta språk.  
Java-program skrivs för det mesta i Java-utvecklingsmiljö och kompileras sedan till "byte-kod".  
Då skapas en .class-fil, som sedan kan infogas som "Java Applet" på t.ex. HTML-sidor.  
Webbläsare som kan tolka Java-program kan utvärdera koden utan att du behöver dekomprimera arkiven.  
Webbläsaren vet då hur detta kommando ska utföras på klientdatorn.  
Ett Java-program kan köras på alla datorer som har en Java-tolk eller -kompilator - t ex en Java-aktiverad webbläsare - oberoende av processortyp och operativsystem.  
Ofta förväxlas JavaScript och Java Applets.  
JavaScript är ett enkelt litet skriptspråk för webbläsare och används t.ex. för visning av rullande text.  
Det beskriver objekt på ett sätt som liknar Java-språket och gör det möjligt för användaren att utsmycka sina HTML-sidor utan att behöva lära sig Java.  
Java Applets är däremot "riktiga" program, som föreligger i form av "Byte Code "enligt beskrivningen ovan.  
Plug-in  
Som plugins (ung.insticksprogram) betecknas sådana utvidgningar av en webbläsare som erbjuder tilläggsfunktioner.  
Mer om plug-ins.  
Plug-in (utförlig förklaring)  
Plug-in är en term som används i olika betydelser.  
Plug-ins i %PRODUCTNAME  
I %PRODUCTNAME ser du gång på gång att objektlister och innehållet på formatmenyerna ändras allt efter situationen.  
Du hittar dem även när du arbetar med rena diagramdokument.  
I det här fallet säger vi att ett diagramdokument körs som plug-in i textdokumentet.  
Ännu tydligare ser du det här funktionssättet om du t.ex. infogar ett textdokument i ett presentationsdokument med Infoga - Objekt - Plug-in.  
Då visas i dokumentfönstret för presentationsdokumentet ett textdokument, och symbollisterna anpassas efter det.  
Plug-ins för programtillägg  
Plug-in-program är i allmänt språkbruk även programtillägg till vissa tillämpningar, som på så sätt utökas med ytterligare funktioner.  
Ofta tillhandahålls import - och exportfilter för olika filformat i form av plug-ins i en plug-in-katalog.  
Även utvidgningar av webbläsaren Navigator från Netscape Communication Corporation kallas plug-in.  
Här rör det sig om externa program, främst på multimedialområdet, som kommunicerar med webbläsaren via ett standardiserat gränssnitt och som också kan läggas in i %PRODUCTNAME -dokument.  
%PRODUCTNAME stöder 32-bitars plug-in-program som kan köras med Netscape Navigator.  
De 32-bitars plug-ins som du har installerat i ett Netscape som finns i ditt system känns automatiskt igen av %PRODUCTNAME och visas i dialogrutan Öppna under Filtyp.  
Om du vill installera 32-bitars plug-ins direkt i %PRODUCTNAME går det att göra med de flesta installationsprogrammen för plug-ins.  
Ange mappen {installpath} / share / plugin som mål, som du skapar och registrerar under Verktyg - Alternativ... - %PRODUCTNAME - Sökvägar.  
Somliga plug-ins kräver dock att Netscape är installerat för att du ska kunna installera dem.  
Proxy  
En proxy är en server i nätverket som fungerar som ett slags cache-minne för dataöverföringen.  
Om du t.ex. kopplar upp dig till Internet från ett företagsnät, sker det vanligen via en proxyserver.  
Webbsidor som tidigare har använts på företaget kan finnas i proxyserverns cache-minne och visas då mycket snabbt på din dator.  
Allt som i så fall måste kontrolleras är om sidan på Internet har uppdateras sedan den sparades senast på proxyservern.  
Om den sida som visas är den aktuella, behöver du alltså inte vänta på att den laddas via en långsam Internet-förbindelse.  
Server  
Servern ställer data, program o.s.v. till förfogande för andra datorer.  
Det finns t.ex. filservrar i lokala nätverk, Internetservrar eller speciella FTP-, e-post - och nyhetsservrar.  
Dessutom kallas även en tillämpning som tillhandahåller data för andra program (klienter) för (application -)server. %PRODUCTNAME Application Server är ett program som körs på en nätverksserver (dator) och som levererar data till %PRODUCTNAME remote-klienter på arbetsstationer.  
SGML  
SGML står för Standard Generalized Markup Language, alltså ungefär "standardiserat allmänt beskrivningsspråk".  
Detta är oberoende av hur dokumenten ser ut senare.  
Ett visst stycke kodas t.ex. som överskrift av första ordningen och efter den ska ett stycke med kodningen bodytext komma.  
SGML definierar vidare hur icke-textinformation, t.ex. videos eller mätvärden, ska överföras till texterna.  
I strukturerade texter kan SGML inte bara definiera strukturen (i DTD = Document Type Definition), utan även kontrollera att den används.  
HTML är en specialtillämpning av SGML.  
Som en följd av detta stöder de flesta webbläsare bara en delmängd av SGML-standarden, samtidigt som alla system som stöder SGML också kan användas för att skapa HTML-sidor.  
De första raderna i ett HTML-dokument innehåller vanligen en SGML-anvisning, som anger att alla följande rader hör till delmängden HTML:  
<!DOCTYPE HTML PUBLIC "- / /W3C / /DTD HTML 3.2 / /EN ">  
SMTP / POP3  
SMTP och POP3 är två mycket använda protokoll för överföring av e-post.  
SMTP (Simple Mail Transfer Protocol) är det vanligaste protokollet med vilket en dator tar kontakt med en e-postserver hos Internetleverantören via modem eller ISDN och överför e-post.  
POP3 (Post Office Protocol, version 3) är ett protokoll som datorn kan använda för att hämta e-post hos Internet-leverantörens e-postserver.  
Style sheets (CSS1 / CSS2)  
Style sheets ("stilmallar") är en nytillkommen funktion i HTML 3-formatet för webbdokument.  
Du kan följa vidareutvecklingen av style sheets på http: / /www.w3.org / Style / Activity.  
Med stilmallar kan du se till att överföringen av formateringen i dina %PRODUCTNAME -dokument fungerar bättre än med de vanliga format taggarna i HTML.  
I stilmallarna finns information om de teckensnitt, teckenstorlekar, radavstånd o.s.v. som ska användas för de olika logiska strukturelementen.  
Detta görs i HTML-koden mellan de nya taggarna <style> och < / style> i form av en lång kommentar.  
I webbläsare som inte stöder stilmallar hoppas det här avsnittet helt enkelt över, medan modernare webbläsare kan utvärdera det.  
Mer om stilar.  
Stilar (ytterligare förklaring)  
Förutom den här typen av infogade (inbäddade) stilmallar kan du göra egna stilmallsfiler, som dina HTML-dokument kan hänvisa till.  
På så sätt kan du bland annat göra stiländringar som är dokumentövergripande genom att ändra i en enda fil.  
CSS (cascading style sheets) är stilmallar som bygger på varandra.  
Sådana stilmallar som är hierarkist ordnade under en huvudstilmall, "ärver" alla attribut hos överordnade mallar och lägger till egna attribut.  
Med hjälp av dynamic HTML kan du lagra objekt ovanpå varandra i tre dimensioner.  
På så vis har du tillgång till bl.a. relativ och absolut placering av sidelement och en synlighet (visibility) som ny egenskap.  
Det finns en omfattande beskrivning på http: / /www.w3.org / pub / WWW / TR / WD-positioning.  
Sökmotor (search engine)  
En sökmotor är en tjänst på Internet som baserar på ett program med vars hjälp du kan söka igenom den oöverskådliga mängden av data på Internet.  
Tags  
HTML -sidor som består av 7-bitars ASCII -text innehåller vissa struktur - och formatanvisningar som kallas taggar.  
De består av nyckelord som är inneslutna av vinkelparenteser och definierade i sidbeskrivningsspråket HTML.  
Många taggar (eng.tags) omfattar en text eller en hyperlänk och utgörs då av en start - och en stopptagg.  
Överskrifter markeras t.ex. med taggen <h1> i början och taggen < / h1> i slutet av överskriftstexten.  
Vissa taggar förekommer inte parvis; t.ex. <br> som anger radbrytning och <img ...> som anger infogning av ett grafikobjekt.  
TCP / IP  
TCP / IP står för Transmission Control Protocol / Internet Protocol.  
TCP är till för upp - och nedkoppling av anslutningar mellan alla datorer i ett nätverk.  
Det styr dataflödet på nätet och ombesörjer en fullständig dataöverföring.  
IP sköter organisation och adressering av data.  
För överföringen delas informationen upp i paket, som sedan sammanfogas hos mottagaren.  
Det här protokollet används både i lokala nätverk och på Internet.  
URL  
En URL (Uniform Resource Locator) anger adressen till ett dokument eller en server på Internet.  
Den allmänna strukturen på en URL varierar beroende på typen men har allmänt formen tjänst: / /värddatornamn:port / sökväg / sida#märke, men alla element behöver inte finnas med.  
En URL kan bland annat vara en FTP-, WWW - (HTTP -), fil - eller e-postadress.  
Web server  
En webbserver är en dator som är ansluten till Internet med ett program som kan visa WWW-dokument och / eller förbereda filer för nedladdning.  
XML  
XML, Extensible Markup Language (utvidgningsbart sidbeskrivningsspråk) är en språkstandard för dokument, utvecklad under ledning av Sun Microsystems.  
Målen för XML var bland andra att XML-dokument utan problem ska kunna användas på Internet och kunna användas av ett stort antal program och vara kompatibla med SGML.  
En utförlig beskrivning av XML finns på http: / /www.w3.org / TR / REC-xml, och på http: / /www.ucc.ie / xml / finns en FAQ-lista.  
Omräkning av måttenheter  
Millimeter  
1 mm = 0,03937008 tum  
1 mm = 0,2362205 pica  
1 mm = 0,1 cm  
1 mm = 56,7 twips  
Pica  
1 pica = 4,233333 mm  
1 pica = 0,4233333 cm  
1 pica = 0,1666667 tum  
1 pica = 12 punkter  
1 pica = 240,029811 twips  
Centimeter  
1 cm = 10 mm  
1 cm = 0,3937008 tum  
1 cm = 2,362205 pica  
1 cm = 28,34646 punkter  
1 cm = 567 twips  
Punkt  
1 punkt = 0,3527778 mm  
1 punkt = 0,03527778 cm  
1 punkt = 0,01388889 tum  
1 punkt = 0,08333333 pica  
1 punkt = 20,00250126 twips  
Tum  
1 tum = 25,4 mm  
1 tum = 2,54 cm  
1 tum = 6 pica  
1 tum = 72 punkter  
1 tum = 1440,18 twips  
Twips  
1 twip = 0,001763668 cm  
1 twip = 0,017636684 mm  
Så hittar du den här funktionen...  
Närliggande ämnen  
Teckenfärg  
Teckenfärg (%PRODUCTNAME Writer)  
Radavstånd:  
1  
Radavstånd:  
1,5  
Radavstånd:  
2  
Upphöjt  
Nedsänkt  
Linjestil  
Linjefärg  
Linjebredd  
Ytstil  
Ytfyllning  
Justera uppe  
Justera nere  
Justera vertikalt i mitten  
Lägg till  
Ta bort  
Ändra kommentar  
Överordnad mapp  
Skapa ny katalog  
Upp en nivå  
Skapa ny mapp  
Standardmapp  
Hopp till föregående anteckning.  
Hopp till nästa anteckning.  
Ladda  
Spara  
Förklaringar av facktermer - Allmän ordlista  
För att det ska bli lättare för dig att komma igång med %PRODUCTNAME, innehåller den här ordlistan förklaringar av de viktigaste facktermerna som du kommer att stöta på.  
Om du precis har börjat arbeta med %PRODUCTNAME stöter du kanske på många obekanta facktermer:  
ODBC, register, SQL och allt möjligt annat.  
I så fall får du reda på det du behöver här.  
Klicka på en av termerna nedan eller bläddra i ordlistan.  
Adabas, ADO, aktivitet, ASCII, Bézierobjekt, bit, bitmap, bågmått (radianer), dBase, DDE, formatering (direkt och indirekt), förankra, grafik, JDBC, kerning, länk, markera, MetaFile, måttenheter (metrik), Native-drivrutin, objekt, ODBC, OLAP, OLE, OpenGL, PNG, primärnyckel, register, relationsdatabas, rotationsfält, RTF, snabbmeny, spara, relativt och absolut, SQL, SQL-severdatabas, %PRODUCTNAME API, talsystem, TWAIN, Unicode, utrullningslist, änkor och horungar.  
Adabas  
Adabas D, version 11, är databasformatet för %PRODUCTNAME -databaser med Windows, Linux och Solaris Sparc.  
Närmare information om Adabas, ytterligare hjälpfiler samt möjligheter att beställa senare versioner finns hos tillverkaren på adressen http: / /www.adabas.com.  
ADO  
Förankra  
Somliga fönster i %PRODUCTNAME kan förankras, t.ex. Stylist, Navigator och Gallery.  
Vid varje kant kan du förankra flera fönster över eller bredvid varandra.  
Du kan ändra den plats som varje förankrat fönster upptar genom att flytta kantlinjerna.  
När du vill ta bort förankringen och förankra igen dubbelklickar du i fönstret och håller ner Kommando Ctrl -tangenten.  
Dubbelklicka på det här sättet på ett tomt område i fönstret.  
I Stylist dubbelklickar du på ett grått ställe i fönstret, t.ex. bredvid ikonerna.  
Det finns det några andra användningstips för hantering av förankringsbara fönster.  
Förankra (utförlig förklaring)  
Vid varje fönsterkant med förankrade fönster finns det två kommandoknappar med vilka du kan visa / dölja eller fixera fönstren.  
Om du använder pilknappen i fönsterkanten för att visa fönstret, visas det tills du döljer det igen med samma knapp.  
Om du visar fönstret genom att klicka på fönsterkanten, aktiverar du funktionen AutoHide.  
Det döljs då automatiskt igen.  
Ta tag i ett fönster i titellisten eller i ett fritt område och flytta fönstret över bildskärmen.  
Om du håller ner Kommando Ctrl -tangenten när du flyttar fönstret, kan fönstret förankras vid kanterna.  
Om du vill förankra ytterligare ett fönster till ett som redan är förankrat, kan du göra det bredvid, ovanför eller under det.  
Lägg märke till hur fönsterkanten ändras.  
Ändringen visar var och med vilken storlek fönstret kommer att förankras.  
Om ett fönster är förankrat kan du göra det till ett fritt fönster igen genom att hålla ner Kommando Ctrl -tangenten och dubbelklicka i ett fritt område.  
ASCII  
Förkortning av American Standard Code for Information Interchange.  
ASCII är en teckenuppsättning för tecken i persondatorer.  
Den består av 128 tecken med bokstäver, siffror, specialtecken och skiljetecken.  
Den utvidgade ASCII-uppsättningen består av 256 tecken.  
Till varje tecken hör ett entydigt nummer som man kallar ASCII-kod.  
På HTML-sidor bör bara tecken från den 7-bitarskodade ASCII-uppsättningen finnas.  
För andra tecken, som t.ex. å, ä, ö, används omskrivningar.  
Så skrivs lilla "ä" som "ä ".  
Exportfiltret i %PRODUCTNAME utför sådana omvandlingar automatiskt.  
Bézier-objekt  
Senare kom sådana kurvor att uppkallas efter honom.  
Med hjälp av kontrollpunkterna och punkterna på kurvan är det lätt att ändra dem med musen.  
Bit  
Bit är en förkortning av "binary digit".  
Detta är den minsta informationsenheten i det binära talsystemet.  
Inom datatekniken sammanförs i många sammanhang 8 bitar till en byte, som behandlas som en enhet.  
Bitmap  
Med bitmap avser man egentligen ett mönster av så kallade bitar.  
I allmänhet menar man ett rastergrafikobjekt eller ett pixelgrafikobjekt.  
Ett sådant objekt är en bild som består av punkter, pixlar, som kan styras oberoende av varandra.  
Vanliga bitmapfilformat är BMP, GIF, JPEG.  
Bågmått  
En vinkel är ett mått på skillnaden i lutning mellan två räta linjer som utgår från samma punkt.  
När man mäter en vinkel utgår man i praktiken från ett helt varv (de räta linjerna sammanfaller) och delar upp den i 360 grader.  
Vid vinkelmätning i bågmått tilldelas varje vinkel en båglängd i "enhetscirkeln"; enheten (som vanligen inte utskrivs) är radian.  
Enhetscirkeln är en cirkel med radien r=1.  
Omkretsen på en cirkel är 2*p*r och för enhetscirkeln är den alltså lika med 2p. (p - "pi "- är en matematisk konstant med det ungefärliga värdet 3,14159265.) Härav gäller följande samband:  
1 grad motsvarar 2*p / 360 = p / 180  
Vinkeln i radianer = gradtalet*p / 180  
Vinkeln i grader = radiantalet*180 / p  
När du använder trigonometriska funktioner måste du tänka på att alla värden beräknas i radianer.  
Eftersom p radianer motsvarar 180 grader, omvandlas gradtalsmått till radianer genom multiplicering med p / 180.  
Omvänt omvandlas radianer till grader genom multiplikation med 180 / p.  
dBase  
Förkortning för Data Base.  
Ett vanligt förekommande databas - och filformat.  
DDE  
DDE står för "Dynamic Data Exchange", alltså dynamiskt datautbyte.  
DDE kan ses som en föregångare till OLE, "Object Linking and Embedding".  
Vid DDE infogas ett objekt i en fil enbart som referens och blir inte "inbäddat".  
En DDE-länk skapas t.ex. när du markerar celler i en %PRODUCTNAME Calc-tabell, kopierar dem till urklippet, sedan byter till ett annat %PRODUCTNAME Calc-dokument och där väljer kommandot Redigera - Klistra in innehåll.  
Markera alternativet DDE-länka i dialogrutan, så infogas cellerna som DDE-länk.  
Varje gång länken aktualiseras, uppdateras det infogade cellområdet genom att cellernas data läses in från ursprungsfilen.  
Formatering  
Med formatering menar man i det här sammanhanget den optiska utformningen av text med ett ordbehandlings - eller designprogram.  
I formateringen ingår bl.a. definition av pappersformat, marginaler, teckensnitt, teckeneffekter, indrag och radavstånd.  
Eftersom det är tidsödande och omständligt att formatera längre texter, finns det i många program - och även i det här %PRODUCTNAME -programmet - särskilda formatmallar.  
Med hjälp av dem kan du formatera ett dokument betydligt snabbare.  
Mer information om direkta och indirekta formateringar.  
Direkta och indirekta formateringar  
Om du formaterar ett dokument utan hjälp av formatmallar, talar man om direkt eller "hård" formatering.  
Med det menar man att texter eller andra objekt - t.ex. ramar eller tabeller - ändras genom att de tilldelas olika attribut.  
Formateringen gäller bara för det markerade området, och alla ändringar måste redigeras var för sig.  
Indirekta eller "mjuka" formateringar gör du däremot inte i själva texten utan genom att tilldela formatmallar.  
Den stora fördelen med det är att du genom att ändra en formatmall ändrar alla objekt (stycken, ramar o.s.v.) som tilldelats den här formatmallen.  
Du kan ta bort direkta formateringar från ett dokument genom att markera allt med tangentkombinationen Kommando Ctrl +A och sedan välja menykommandot Format - Standard.  
Grafik, vektorgrafik och pixelgrafik  
I datorvärlden skiljer man mellan vektorgrafik och pixelgrafik.  
Bilder med vektorgrafik består av anvisningar såsom "dra en linje med färgstyrka A och färg B från punkten med koordinaterna (C,D) till punkten (E,F)".  
Sådana bilder är oberoende av bildskärmsupplösningen, vilket betyder att de alltid har samma kvalitet (inom ramen för utmatningsmediets prestanda) oavsett förstorings - eller förminskningsgrad.  
I %PRODUCTNAME skapar du vektorgrafikobjekt via Arkiv - Nytt - Presentation respektive Teckning.  
Bilder med pixelgrafik består av intilliggande pixlar, bildpunkter, som kan ha olika färger.  
Sådana bilder har alltid definierade mått, t ex 800 pixlar bred och 600 pixlar hög, varvid en pixel är den minsta måttenheten.  
När man förstorar pixelgrafikobjekt, i exemplet till låt säga 1000 x 800, uppstår problem.  
Man kan inte bara förstora varje enskild pixel, eftersom den har en given storlek som beror av utmatningsmediet (t ex bildskärmen).  
Alltså måste man dubblera vissa pixlar men inte andra, och eventuellt även beräkna övergångsfärger.  
Den processen gör att kvaliteten blir lidande.  
Ändå är användningen av pixelgrafik mycket vanlig, eftersom kameror, skannrar och liknande utrustning skapar pixelgrafik.  
Program för retuschering av pixelgrafik finns på alla möjliga kvalitets - och prisnivåer.  
Du skapar pixelgrafik i %PRODUCTNAME Draw genom att välja kommandot Arkiv - Exportera och sedan ett motsvarande filformat, t.ex. JPG.  
JDBC  
JDBC står för Java DataBase Connectivity och är precis som ODBC ett protokoll för åtkomst av databassystem.  
Skillnaden mot ODBC är bara att drivrutinen för JDBC är programmerad i Java och därmed plattformsoberoende.  
Kerning  
Kerning är en engelsk beteckning för att minska eller öka avståndet mellan bokstavspar, t.ex. mellan V och a.  
På så sätt uppnår man en optisk utjämning av teckenbilden.  
Kerningtabellerna innehåller information om för vilka bokstavspar avståndet ökas eller minskas och hur mycket.  
De här tabellerna är i allmänhet en del av definitionen av ett teckensnittet.  
Metafil  
Windows Metafile Format (WMF) är ett grafikformat som har utvecklats för Microsoft Windows.  
WMF-grafikfiler kan innehålla både bitmap - och vektordata.  
I %PRODUCTNAME Draw och %PRODUCTNAME Impress används metafilformatet som vektorformat.  
Native-drivrutin  
%PRODUCTNAME innehåller s.k. native-drivrutiner för speciella databassystem.  
Med hjälp av en native-drivrutin får du som användare direkt åtkomst till respektive databasklient.  
Objekt  
Ett objekt är ett element på bildskärmen som innehåller information.  
Det kan t.ex. röra sig om användningsdata som text eller grafik.  
Objekt är självständiga och påverkar inte varandra.  
Det finns särskilda kommandon för varje objekt som innehåller data.  
Ett grafikobjekt förses t.ex. med kommandon för bildredigering och en tabell med kommandon för beräkning.  
ODBC  
ODBC står för Open DataBase Connectivity, d.v.s. ungefär öppen databasanslutning.  
Detta är ett standardiserat protokoll, med vars hjälp tillämpningsprogram kommer åt databassystem.  
Som frågespråk används SQL (Structured Query Language = språk för strukturerade frågor).  
Den översätts i så fall till SQL av %PRODUCTNAME.  
De nödvändiga 32-bitars ODBC-funktionerna installerar du i operativsystemet med hjälp av ett setup-program från databastillverkaren.  
Egenskaperna ställer du in på kontrollpanelen.  
OLAP  
OLAP är en förkortning av O n l ine A nalytical P rocessing, d.v.s. analytisk onlineredigering.  
Det rör sig om särskilda program för dataanalys i databaser.  
Med OLAP-program kan du analysera olika dimensioner i flerdimensionella datastrukturer, t.ex. göra trendanalyser.  
Huvudkomponenten i OLAP är OLAP-servern, som befinner sig mellan klienten och databashanteringssystemet (DBMS; Database Management System).  
OLAP-servern förstår hur data i en databas är organiserade och förfogar över särskilda funktioner för analys av dessa data.  
Det finns OLAP-servrar för nästan alla databassystem.  
OLE  
Förkortning av Object Linking and Embedding (länkning och inbäddning av objekt).  
Objekt kan länkas till ett måldokument eller om så önskas "bäddas in" där.  
Vid inbäddning infogas en kopia av objektet i måldokumentet tillsammans med uppgifter om källprogrammet.  
Det gör att källprogrammet öppnas om du dubbelklickar på objektet, och på så vis kan du komma åt att redigera det.  
OpenGL  
OpenGL är ett språk för 3D-grafik, ursprungligen utvecklat av SGI (Silicon Graphics Inc.).  
Det finns två mycket spridda tillämpningar av OpenGL, nämligen Microsoft OpenGL, utvecklat för Windows NT, och Cosmo OpenGL från SGI.  
Det senare är ett plattformsoberoende grafikspråk för alla datorer, även sådana som inte har någon särskild maskinvara för 3D-grafik.  
PNG  
PNG (uttalas "Ping") står för Portable Network Graphics.  
Det är ett dataformat för lagring av pixelgrafik vars betydelse på Internet sakta med säkert växer.  
Grafikobjekten komprimeras med en valfri faktor, men i motsats till JPG-formatet sker komprimeringen alltid utan förlust av bilddata.  
PNG kan lagra 24 - och 8-bitars färgbilder, gråskalor och svartvita bilder; om så önskas med alfakanaler för transparensinformation.  
Vid överföring av PNG-bilder med egenskapen "interlaced" visas till att börja med var n:te bildlinje eller -kolumn, och efterhand fylls luckorna ut.  
Primärnyckel  
En primärnyckel är till för entydig identifiering av ett databasfält.  
Denna entydiga identifiering av databasfält används i relationsdatabaser, där identifieringen av data i den ena tabellen kan användas för åtkomst av data i en annan.  
Om en annan tabell innehåller en referens till en primärnyckel, betecknar man den referensen som sekundärnyckel.  
I %PRODUCTNAME definierar du primärnycklar i utkastvyn av en tabell genom att välja motsvarande kommando för det markerade fältet på snabbmenyn till ett radhuvud.  
Relationsdatabas  
Relational Database Management System) är ett databassystem där data hanteras i form av tabeller som är kopplade till varandra.  
En väl planerad databas kan vara uppbyggd så att varje uppgift bara behöver matas in en gång men ändå kan granskas i flera olika sammanhang.  
Ett klassiskt exempel på en relationsdatabas är tabeller med kunddata, varudata och fakturadata relaterade till beställningar.  
Bokföringstabellen innehåller inte namnen på kunder och varor utan hänvisningar till motsvarande dataposter i andra tabeller.  
Länkningen görs via gemensamma datafält med t ex kundnummer och artikelnummer.  
Register  
Register är en typografisk term.  
Med det menas att raderna på den ena sidan på bladen i böcker, tidskrifter osv har exakt samma position som motsvarande rad på den andra sidan.  
På det viset undviker man att det uppstår grå fält mellan raderna (på grund av att raderna på baksidan svagt skiner igenom), vilket försvårar läsningen.  
Man talar även om register när alla rader som ligger bredvid varandra i textspalter har samma höjd. (Ett annat och kanske vanligare uttryck är att raderna linjerar med varandra.)  
Om du ställer in registret för stycken, sidor eller stycke - resp. sidformatmallar i ett textdokument justeras radernas baslinjer så att de passar in i det vertikala radrastret i styckeformatmallen som du har angett som referensmall.  
Baslinjerna för intilliggande rader i alla stycken med register är fortfarande justerade på samma höjd (de linjerar).  
RTF  
Förkortning av Rich Text Format ("fylligt "textformat).  
Filformat avsett för tillämpnings - och plattformsoberoende utbyte av formaterade textdata.  
En speciell egenskap är att formateringarna ger direkt läsbar textinformation.  
Filstorleken är naturligtvis betydligt större än för rent ASCII-format (som också det är tillämpnings - och plattformsoberoende).  
Änkor och horungar  
Änkor och horungar är typografiska beteckningar av mycket gammalt datum.  
En horunge är när sista raden i ett stycke står överst på nästa sida.  
I ett textdokument i %PRODUCTNAME kan du undvika dessa fenomen automatiskt genom att ställa in styckeformatmallen på det sättet.  
Du kan t.o.m. välja hur många rader som minst måste förekomma tillsammans på en sida.  
Markera  
Nästan alla kommandon i %PRODUCTNAME, t.ex. för formatering av text n %PRODUCTNAME Writer, refererar till markering.  
Text markerar du t.ex. med musen genom att hålla ner musknappen och stryka över texten.  
Den markerade texten visas inverterad.  
Spara relativt och absolut  
I olika dialogrutor (t.ex. Redigera - AutoText) kan du välja om du ska spara filer relativt eller absolut.  
När du väljer bör du ta hänsyn till hur dokumenten i fråga ska användas.  
Mer information om att spara relativt och absolut.  
Spara relativt och absolut  
Om du väljer att spara relativt, kommer referenserna till inbäddade grafikobjekt eller andra filbaserade objekt i dokumentet att infogas i en form som utgår från dokumentets plats i filstrukturen.  
Det spelar ingen roll om den filstrukturen befinner sig på t.ex. enhet C: eller enhet D: respektive volym HD1, HD2 eller någon annanstans.  
Filerna kommer hur som helst att hittas (så länge referensfilen finns kvar i samma enhet eller volym).  
Detta är särskilt viktigt om du lägger upp en filstruktur på en Internet-server, t.ex. i en hemsidesmapp hos Internet-leverantören.  
Om du föredrar att spara absolut, blir alla referenser till andra filer absoluta, d.v.s. de utgår från respektive enhet, volym eller rotkatalog.  
Det har fördelen att du kan flytta dokumentet där referenserna finns till andra kataloger eller mappar på datorn utan att referenserna blir ogiltiga.  
Det är å andra sidan bättre att referenser sparas relativt i stället för absolut för dokument som ska vara tillgängliga på en annan dator, som kan ha en helt annan katalogstruktur och andra enhets - eller volymbeteckningar.  
SQL  
"Structured Query Language" är ett strukturerat frågespråk för databaser.  
I %PRODUCTNAME kan Du formulera Dina frågor till databasen som Du vill, antingen med SQL eller med musen.  
SQL-databas / SQL-server  
En SQL-databas är ett databassystem som tillhandahåller ett SQL -gränssnitt.  
Därför betecknar man dem även SQL-serverdatabaser eller kort och gott SQL-servrar.  
I %PRODUCTNAME kan du integrera externa SQL-databaser.  
De kan finnas antingen på hårddisken eller i nätverket.  
Åtkomsten sker antingen via ODBC eller via en native-drivrutin integrerad i %PRODUCTNAME.  
%PRODUCTNAME API  
%PRODUCTNAME API (Application Program Interface) är gränssnittet för programmering av %PRODUCTNAME.  
Den ger programstyrd åtkomst till alla delar av %PRODUCTNAME och möjliggör utveckling av egna tilläggsmoduler. %PRODUCTNAME API kan nås både från Java och från Microsofts Component Object Model.  
Aktivitet  
Aktivitet (eng. task) är den allmänna beteckningen på en begränsad del av ett programs funktioner och åtgärder.  
Ur operativsystemets perspektiv är bl.a. de program som just körs aktiviteter; för ett program som %PRODUCTNAME är bl.a. de enskilda dokumenten aktiviteter.  
I en möteskalender kan de införda uppgifterna betecknas som aktiviteter.  
TWAIN  
TWAIN är ett standardiserat protokoll och gränssnitt för tillämpningsprogram (API) för kommunikation mellan enheter som bearbetar bilder (skannrar, digitalkameror) och programvaran.  
TWAIN stöds för närvarande bara av Windows.  
Se http: / /www.mostang.com / sane /.  
Unicode  
Unicode är ett system där tecken och element från alla kända skrivkulturer och teckensystem har förts samman.  
Varje tecken eller element kodas till ett tal som är två byte långt.  
Genom UTF-16 Extension kan över en miljon olika tecken återges.  
De relativt trånga gränserna för enskilda teckenuppsättningar hör därmed till det förgångna.  
Med Unicode kan olika språk blandas utan problem.  
Det finns mer information på Unicode-konsortiets hemsida: http: / /www.unicode.org.  
Länk  
Det är bara tillgängligt när det finns minst en länk i det aktuella dokumentet.  
Ett objekt, t.ex. ett grafikobjekt, som du infogar i dokumentet kan antingen kopieras dit eller infogas som länk.  
Vid direkt kopiering ökar dokumentfilens omfång med minst objektets storlek.  
Du kan spara dokumentet och öppna det på en annan dator, och det infogade objektet finns fortfarande på sin plats.  
Om du infogar objektet som länk, skapas bara en referens till filnamnet.  
Dokumentets filstorlek ökar bara med det utrymme som länken upptar.  
Men om du öppnar dokumentet på en annan dator, måste den länkade filen finnas på exakt den adress som referensen anger för att objektet ska kunna visas.  
I dialogrutan Redigera länkar kan du se vilka filer som är länkade till dokumentet.  
Du kan även radera länkarna här om du vill.  
Talsystem  
Ett visst talsystem kännetecknas av det antal siffertecken som står till förfogande för skrivning av tal.  
Detta antal siffertecken är den matematiska basen för talsystemet.  
Det system som vi använder till vardags är decimalsystemet, som har basen 10 och tio siffertecken (0-9).  
Vidare har vi i binärsystemet med basen 2 (siffrorna 0 och 1) och hexadecimalsystemet med basen 16 (siffrorna 0-9 och bokstäverna A-F) två viktiga talsystem.  
Namn på lister  
Ikon på verktygslisten:  
Ikon på textobjektlisten:  
Ikon på objektlisten:  
Ikon på objektlisten i diabildsvyn:  
I %PRODUCTNAME är det lätt att ändra menyer, ikoner och symbollister.  
Om du drar nytta av den möjligheten avviker din konfiguration från den som beskrivs här.  
Asiatiska specialfunktioner  
De här kommandona visas bara om du har aktiverat stödet för asiatiska språk under Verktyg - Alternativ - Språkinställningar - Språk.  
Snabbmenyer  
Klipp ut  
Klipper ut det markerade objektet och placerar det i urklippet.  
Därifrån kan det infogas med Klistra in.  
Klistra in  
Infogar det element som du kopierat till urklippet med Kopiera.  
Du kan bara välja det här kommandot när det är någon mening att infoga innehållet i urklippet vid infogningspositionen.  
Lägg till...  
Öppnar en undermeny i Gallery där du kan välja bland alternativen Kopia och Länk.  
När du har valt ett av alternativen i undermenyn kopieras det markerade grafikobjektet till det aktuella dokumentet eller så skapas en länk i dokumentet.  
Om någonting är markerat i ditt dokument, t.ex. det senast inklistrade grafikobjektet, ersätts som vanligt det markerade objektet vid en ny inklistring.  
Bakgrund  
Med denna funktion infogar du det markerade grafikobjektet som bakgrundsbild.  
Med undermenyalternativen Sida och Stycke bestämmer du om grafikobjektet ska ligga i bakgrunden på hela sidan eller bara bakom det aktuella stycket.  
Kopiera  
Kopierar det markerade elementet till urklippet.  
Radera  
Raderar den aktuella markeringen.  
Vid en multipel markering raderas samtliga markerade objekt.  
Innan raderingen får du en kontrollfråga.  
Beroende på sammanhanget raderas objektet fysiskt från datamediet eller också tas det bara bort från visningen av objektet.  
Om du väljer kommandot Radera i Gallerys tas posten bort från visningen i Gallery, men filen rörs inte.  
Sökning...  
Öppnar en undermeny där du kan välja om du vill skapa sökningen i utkastläge eller med hjälp av AutoPiloten  
Formulär  
Öppnar en dialogruta där Du kan välja typ av formulär.  
Tabell  
Öppnar en undermeny där Du kan välja om Du vill skapa tabellen i utkastläge eller med hjälp av AutoPiloten.  
Tabellvisning  
Här kan Du öppna ett fönster för att definiera en ny vy över en tabell som Du t ex har åtkomst till via en databasserver.  
Öppna  
Med det här kommandot öppnar du det markerade objektet i en egen aktivitet.  
%PRODUCTNAME databas (namn: [Kortnamn])  
Här anger Du om databasen ska registreras med ett kort namn eller inte.  
Om databasen är registrerad är kommandot förbockat.  
Ytterligare information finns i hjälpen för %PRODUCTNAME under rubriken Databasnamn.  
Byt namn  
Tillåter att du byter namn på det markerade objektet.  
När du har valt kommandot Byt namn markeras namnet.  
Du kan skriva in ett nytt namn direkt eller placera markören i början eller slutet av namnet med piltangenterna och ta bort eller lägga till delar eller flytta markören till ett annat ställe.  
Uppdatera  
Klicka på den här posten för att uppdatera visningen i det aktuella fönstret eller det markerade fönstret.  
Förhandsvisning  
Det element som är markerat visas i Gallery i maximal storlek.  
Dubbelklicka på förhandsvisningen för att återgå till normalvy i Gallery.  
Skapa länk  
Det här kommandot går att aktivera när ett objekt är markerat.  
Länken får namnet "Länk till xxx" (xxx står för objektets namn).  
Menykommandon  
Kommandona för att till exempel redigera, se, placera, formatera och skriva ut ett dokument eller dokumentets innehåll, går bara att använda om dokumentet är öppet och aktivt.  
Aktivt innebär här att dokumentet måste vara i förgrunden på bildskärmen.  
Om du vill använda kommandon till ett objekt i dokumentet måste objektet vara markerat.  
Det betyder att alltid de menykommandon står till förfogande som är relevanta i respektive sammanhang.  
Om till exempel ett grafikobjekt är markerat i dokumentet, hittar du alla menykommandon som används till att redigera grafik.  
Du ser alltid bara de menyposter som går att använda.  
De andra inaktiva menyposterna är dolda.  
Om du vill se de inaktiva menykommandona i grått kan du välja Verktyg - Alternativ - %PRODUCTNAME - Vy och markera rutan Inaktiva menyposter.  
Information om import - och exportfilter  
I %PRODUCTNAME kan du inte bara öppna och skriva i de egna XML-formaten utan även i många externa format.  
Under UNIX kan en del filformat inte identifieras automatiskt.  
Det kan förekomma situationer när du själv måste välja filtyp i dialogrutan Öppna.  
Anta att du t.ex. har en databastabell i textformat, som du också vill öppna som databastabell.  
I det här fallet väljer du inte bara fil utan även filtypen "".  
Det är bara då som dialogrutan Textimport av en databastabell öppnas.  
Där kan du t.ex. välja alternativet Engelska (US).  
Oberoende av systemspråk försöker nu programmet att tolka innehållet som tal formaterade enligt amerikansk standard.  
De engelska månadsnamnen känns i varje fall igen automatiskt.  
Basic-makron i MS Office-dokument  
Under Verktyg - Alternativ - Ladda / spara - Microsoft Office kan du bestämma vad som ska hända med VBA Makro Codes i MS Office-dokument.  
VBA-makron går inte att köra under %PRODUCTNAME; de måste först konverteras och anpassas.  
Ofta vill du kanske bara ändra det synliga innehållet i en Word-, Excel - eller Power Point-fil med hjälp av %PRODUCTNAME och sedan spara filen i Microsoft Office-format igen, utan att ändra makron som finns i filen.  
Du kan ställa in hur %PRODUCTNAME ska göra:  
Antingen sparas VBA-makrona temporärt i kommenterad form som en subrutin till %PRODUCTNAME och skrivs tillbaka korrekt när dokumentet sparas i MS Office-format, eller så kan du välja att %PRODUCTNAME tar bort makrona vid laddningen.  
Det senare alternativet är naturligtvis ett effektivt skydd mot Virus i Microsoft Office-dokument.  
Anmärkningar kring %PRODUCTNAME :s egna format  
I %PRODUCTNAME Writer kan du fr.o.m. version 5.0 ladda och spara betydligt större textdokument än i tidigare versioner.  
Därför kan ett försök att spara ett mycket stort dokument i ett äldre %PRODUCTNAME Writer-format leda till att ett felmeddelande visas.  
Anmärkningar beträffande externa format och filtyper  
En del filter går att välja i dialogrutorna för att öppna och spara dokument, trots att de inte är installerade.  
När du väljer ett sådant filter får du en upplysning om att du kan installera detta filter i efterhand.  
Om du vill installera fler filter eller ta bort enskilda filter från installationen, avslutar du %PRODUCTNAME och kör setupprogrammet för %PRODUCTNAME %PRODUCTVERSION.  
Då visas en dialogruta där du kan lägga till eller ta bort enskilda komponenter i %PRODUCTNAME.  
Grafikfilter finns under "Valfria komponenter".  
Import och export av textdokument  
Du kan också spara dina egna texter i Word-format.  
Men allt som man kan göra i %PRODUCTNAME Writer kan inte överföras till MS-Word och allt kan inte importeras.  
När du exporterar dispositioner i %PRODUCTNAME Writer till Word-format följer bara den första dispositionen per giltighetsområde i en sidmall med, eftersom Word inte kan bearbeta flera dispositioner.  
Samtliga därpå följande dispositioner får därför samma layout som den första.  
Word kan inte heller använda grafikobjekt som bullets (punkter).  
Motsvarande gäller för tecken före och efter siffror.  
I normala fall går det att importera utan problem.  
Även redigeringsinformation och kontrollfält (controls) importeras (och exporteras), så att nya infogade texter, raderade texter och ändrade teckenattribut i ett Word-dokument kan identifieras av %PRODUCTNAME och ges olika färger beroende på vem som gjort ändringarna.  
Även information om när redigeringarna gjordes följer med vid importen.  
Det kan dock hända att attribut går förlorade.  
Naturligtvis går det även att importera och exportera RTF -filer.  
Syftet med det här filformatet är att man ska kunna flytta formaterade texter mellan olika program och plattformar.  
På så vis kan formateringar överföras mellan de flesta program.  
Med det här formatet arbetar också urklippet när du klistrar in ett område från %PRODUCTNAME Calc i %PRODUCTNAME Writer via DDE.  
Textfiltret Text - kodad används till att öppna och spara textdokument med annan kodning för teckenuppsättningar.  
Filtret har en dialogruta där du kan ställa in teckenuppsättning, standardteckensnitt, språk och styckebrytning.  
Import och export i HTML-format  
När du exporterar inramningar i HTML-dokument, t.ex. en styckeinramning, exporteras linjer som är 1 pixel breda, eftersom Netscape Navigator och MS Internet Explorer inte kan identifiera tunnare linjer.  
Vid en import omvandlas en linje med bredden 1 pixel till en linje med bredden 0,05 pt.  
Med %PRODUCTNAME Writer kan du också infoga fot - och slutnoter i HTML-dokument.  
Fot - och slutnotstecknen exporteras som hyperlänkar.  
För att även okända tecken ska kunna sparas i HTML-dokument används noter.  
Varje not som börjar med "HTML:..." och slutar med "> "behandlas som HTML-kod, men exporteras utan dessa beteckningar.  
Bakom "HTML:..." kan det stå flera taggar och mellan dessa valfri text.  
Omljud konverteras till ANSI-teckenuppsättningen.  
Även vid import läggs det upp anteckningar (t ex för metataggar för vilka det inte finns plats i dokumentinformationen eller okända taggar).  
HTML-importen i %PRODUCTNAME Writer kan läsa filer som finns i UTF-8 - respektive UCS2-teckenkodning.  
Alla tecken som finns i ANSI-teckenuppsättningen eller i systemets teckenuppsättning visas.  
Vid export till HTML används den teckenuppsättning som du väljer under Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet.  
Tecken som inte finns där skrivs i ersättningsformen "Ӓ" som visas korrekt av moderna webbläsare.  
När du exporterar sådana tecken får du en varning om det.  
Om du har ställt in Netscape Navigator 4.0, MS Internet Explorer 4.0 eller %PRODUCTNAME Writer som exportalternativ via Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet, exporteras alla viktiga teckenattribut som direkta attribut (t.ex. textfärg, teckenstorlek, fet, kursiv o.s.v.) i CSS1-styles. (CSS betyder Cascading Style Sheets.  
Även importen följer denna standard.  
Det innebär att Du innan fontstorleken kan ange värden för "font-style" (italic, none), "font-variant "(normal, small-caps) och "font-weight" (normal, bold).  
Om något av värdena inte anges återställs det.  
t ex font: bold italic small-caps 12pt / 200% Arial, Helvetica kopplar om till fet, kursiv, små kapitäler, 12pt-skrift, dubbla radavstånd med fontfamiljen Arial eller Helvetica om Arial inte skulle finnas.  
10pt växlar över till ett 10 punkters teckensnitt som är fetstilt, kursivt och har små kapitäler.  
Om MS Internet Explorer 4.0 eller %PRODUCTNAME Writer ställts in som exportalternativ, exporteras kontrollfältens storlek och dessas avstånd till innehållet som Styles (utskriftsformat).  
När det gäller storlek används CSS1-egenskaperna "width" och "height ".  
Om avstånden inte är lika stora används egenskaperna "margin-left", "margin-right", "margin-top" och "margin-bottom ".  
Avståndet från grafik, PlugIns och Appletprogram till innehållet kan du ställa in individuellt för %PRODUCTNAME Writer och MS Internet Explorer 4.0.  
Om det övre / nedre eller högra / vänstra avståndet har olika inställning, exporteras avstånden i ett "STYLE"-alternativ för respektive tagg som CSS1-egenskaperna "margin-top", "margin-bottom", "margin-left" och "margin-right ".  
Genom användningen av CSS1-utökningar för absolut placerade objekt understöds också textramar.  
Men detta gäller bara för export-webbläsarna Netscape Navigator 4.0, MS Internet Explorer 4.0 och %PRODUCTNAME Writer.  
Textramar som grafik, plug-ins appletprogram och flytande ramar kan justeras, men inte teckenbundna ramar.  
Textramar exporteras som "<SPAN>" - eller "<DIV> "-tag om de inte innehåller några kolumner.  
Om de innehåller kolumner exporteras textramar som "<MULTICOL>".  
Vid HTML-export används den måttenhet som ställts in för CSS1-egenskaper i %PRODUCTNAME.  
Måttenheten kan ställas in separat för text - och HTML-dokument under Verktyg - Alternativ - Textdokument - Allmänt respektive Verktyg - Alternativ - HTML-dokument - Vy.  
Antalet exporterade decimaler beror på enheten:  
Måttenhet  
Namn på måttenheten i CSS1  
Maximalt antal decimaler  
millimeter  
mm  
2  
centimeter  
cm  
2  
tum  
in  
2  
pica  
pc  
2  
punkt  
pt  
1  
Webbsidesfiltret i %PRODUCTNAME stöder en del funktioner i CSS2.  
För att du ska kunna utnyttja dem måste du aktivera export av utskriftslayout under Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet.  
I HTML-dokument kan du då använda formatmallarna "första sida", "vänster sida" och "höger sida ", förutom HTML-sidformatmallen.  
Syftet med de här formatmallarna är att du ska kunna ange olika sidstorlekar och kanter för den första, den vänstra och den högra sidan.  
Import och export av numreringar  
Om du väljer exportalternativet "%PRODUCTNAME Writer" eller "Internet Explorer "under Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet exporteras numreringarnas indrag som "margin-left "-CSS1-egenskaper i STYLE-attributet för <OL> - och <UL>-taggar.  
Egenskapen anger differensen i förhållande till indraget på den direkt ovanförliggande nivån.  
Ett vänsterstyckeindrag exporteras inom numreringar som en "margin-left "-CSS1-egenskap.  
Förstaradsindragningar ignoreras vid numreringar och exporteras därför inte heller.  
Import och export av tabellfiler  
Vid export syns hela formeln och den raderade referensen får en hänvisning till det refererade (#REF).  
På motsvarande sätt skapas vid import en #REF! för referensen.  
Import och export av grafikfiler  
På liknande sätt som för HTML-dokument kan du bestämma om du vill använda ett filter med eller utan tillägget (%PRODUCTNAME Impress) i namnet när du öppnar en %PRODUCTNAME -grafikfil.  
I det andra fallet öppnas filen som ett %PRODUCTNAME Draw-dokument.  
EPS-grafik importeras och förhandsvisas sedan.  
Förhandsvisningen skrivs ut med andra skrivare.  
Vid export av EPS-grafik kan du skapa en förhandsvisning i TIFF - eller EPSI-format.  
Om EPS-grafik exporteras tillsammans med annan grafik i EPS-format integreras filen i den nya filen i oförändrat skick.  
Vid import och export av grafikfiler i TIFF-format tas också hänsyn till s k multipage-tiff.  
Det rör sig i detta fall om en samling enskilda bilder i en enda fil, t ex enskilda sidor från ett fax.  
Vissa alternativ i %PRODUCTNAME Draw och %PRODUCTNAME Impress når du via menyn Arkiv - Exportera.  
PostScript  
Om du vill exportera ett dokument eller ett grafikobjekt i ett PostScript-format gör du så här:  
Om det inte redan gjorts installerar du en drivrutin för PostScript, t.ex. drivrutinen till Apple LaserWriter.  
Skriv ut dokumentet med menykommandot Arkiv - Skriv ut I dialogrutan väljer du PostScript-skivaren och klickar i rutan Skriv ut till fil.  
När du skriver ut skapas nu en PostScript-fil.  
XML-filformat  
Standardfilformatet för att öppna och spara dokument i %PRODUCTNAME är ett XML-filformat.  
Namnen på XML-filformaten  
Om du inte väljer någon annan filtyp i dialogrutorna för att spara och öppna %PRODUCTNAME -dokument, använder %PRODUCTNAME följande XML-filformat:  
Användning  
Filnamnstillägg  
%PRODUCTNAME Writer  
*. sxw  
%PRODUCTNAME Writer-mallar  
*.stw  
%PRODUCTNAME Calc  
*.sxc  
%PRODUCTNAME Calc-mallar  
*.stc  
%PRODUCTNAME Impress  
*.sxi  
%PRODUCTNAME Impress-mallar  
*.sti  
%PRODUCTNAME Draw  
*.sxd  
%PRODUCTNAME Draw-mallar  
*.std  
%PRODUCTNAME Math  
*.sxm  
Samlingsdokument  
*.sxg  
De här filnamnstilläggen gör att det är lättare att skilja många filer med olika filtyper åt i en katalog.  
Dessutom talar beteckningen om att det rör sig om komprimerade XML-filer som först måste dekomprimeras innan t.ex. en textredigerare kan läsa dem.  
Om du vill arbeta permanent med ett annat filformat kan du definiera det som standard.  
Du kanske t.ex. inte vill använda *.sxw-formatet som standard för att öppna och skriva i %PRODUCTNAME Writer utan ett *.doc-format.  
Under Verktyg - Alternativ - Ladda / spara - Allmänt kan du välja alternativa filformat för alla %PRODUCTNAME -dokumenttyper.  
XML-filens struktur  
XML-filformaten i %PRODUCTNAME är komprimerade enligt ZIP-metoden.  
Använd ett valfritt dekomprimeringsprogram för att "packa upp" innehållet i en XML-fil med dess underordnade kataloger.  
En struktur visas som ser ut ungefär så här (se bild).  
Textinnehållet i dokumentet står i content.xml.  
Du kan t.ex. titta på den här filen med en ren textredigerare.  
Standard är att content.xml sparas utan indrag i början av raden så att det inte tar så lång tid att spara och öppna.  
Under Verktyg - Alternativ - Ladda / spara - Allmänt kan du ändra detta så att raderna sparas med indrag.  
Du kan mata in den här informationen under Arkiv - Egenskaper.  
Om du sparar ett dokument krypterat är meta.xml den enda filen som inte krypteras.  
I settings.xml finns det mer information om inställningar för det här dokumentet, t.ex. om skrivaren, om registrering av ändringar, den anslutna datakällan med mera.  
I styles.xml kan du se vilka formatmallar som har definierats för dokumentet.  
Filen meta-inf / manifest.xml beskriver XML-filens struktur.  
Det kan finnas fler filer i ett komprimerat filformat.  
Illustrationer står t.ex. i en underordnad katalog som heter Pictures, Basic-kod i en underordnad katalog som kallas Basic och anslutna Basic-bibliotek finns i andra underordnade kataloger till Basic.  
Definition av XML-formaten  
DTD (Document Type Description)-filerna finns i {installpath} / share / dtd {installpath }\share\dtd.  
Tänk på att formaten är licensbelagda.  
Information om licenserna finns i början av DTD-filerna.  
Detaljerad information finns på OpenOffice.org -webbsidan.  
Installationen av %PRODUCTNAME är ofullständig  
Om den här dialogrutan öppnas automatiskt upptäcktes det vid starten av %PRODUCTNAME att det saknas viktiga filer eller så har de inte registrerats korrekt i systemet och att felet inte kunde avhjälpas automatiskt.  
Försök att åtgärda felet på följande sätt:  
Avsluta %PRODUCTNAME och öppna %PRODUCTNAME Setup.  
Välj alternativet Reparation.  
komponenter som saknas  
I den här listan visas de komponenter som för närvarande saknas eller som inte registrerats korrekt i systemet.  
Gör alltid den här kontrollen vid start av %PRODUCTNAME  
Ta bort markeringen om det inte längre ska göras någon kontroll vid start av %PRODUCTNAME.  
Se även...  
Meny Verktyg - Scenarion  
På hjälpsidan till %PRODUCTNAME allmänt finns modulberoende anvisningar som t.ex. hur du arbetar med fönster och menyer, anpassar %PRODUCTNAME, datakällor, Gallery, dra-och-släpp och så vidare.  
Om du vill ha hjälp till en annan modul så väljer du först ut den här andra modulen i kombinationsfältet i navigationsområdet.  
JPEG-alternativ  
I denna dialogruta gör Du inställningar för export och import av filer i JPEG-format.  
Kvalitet  
Välj önskad grafikkvalitet.  
Kvalitet  
Markera export - respektive importkvaliteten i rotationsfältet.  
Värdet 0 betyder minimal kvalitet och minimal filstorlek, värdet 100 betyder maximal kvalitet och filstorlek.  
Färgupplösning  
Markera önskad färgupplösning.  
Gråskalor  
Välj den här rutan om du vill exportera eller importera grafik i gråskalor.  
True Colors  
Välj den här rutan om du vill behålla originalfärgerna i JPEG-filen vid export respektive import.  
Mer information om filtrering finns i avsnittet om import - och exportfilter.  
SVM / WMF / PICT / MET-alternativ  
Här markerar Du exportalternativ.  
Läge  
I detta område väljer Du läge för filexport.  
Original  
Klicka här om Du vill behålla originalstorleken.  
Storlek  
Markera denna ruta om Du vill ändra storleken.  
Storlek  
Detta område är bara aktivt om Du markerade alternativet Storlek under Läge.  
Bredd  
Ange bredden här.  
Höjd  
Ange höjden här.  
Mer information om filtrering finns i avsnittet om import - och exportfilter.  
Det innehåller följande undermenyer:  
1Bit-tröskelvärde  
Objektet färgläggs i svart och vitt.  
Alla ljusstyrkenivåer under medelvärdet blir svarta och alla över blir vita.  
1Bit-Ditrering  
Objektet färgläggs med ett rutnät av svarta och vita punkter.  
4Bit-gråskalepalett  
Objektet färgläggs med 16 gråskalor motsvarande originalets ljusstyrka.  
4Bit-färgpalett  
Objektet färgläggs med 16 färger som bäst motsvarar originalfärgerna.  
8Bit-gråskalepalett  
Objektet färgläggs med 256 gråskalor motsvarande originalets ljusstyrka.  
8Bit-färgpalett  
Objektet färgläggs med 256 färger som bäst motsvarar originalfärgerna.  
24Bit-TrueColor  
Gör det möjligt att färglägga ett objekt med ett urval av 16 miljoner färger.  
BMP-alternativ  
I denna dialogruta gör Du inställningar för export av filer i BMP-format.  
Färgupplösning  
Här väljer Du färgupplösning.  
Färgupplösning  
I denna listruta hittar Du alla upplösningsalternativ som finns tillgängliga.  
RLE-kodning  
Klicka här om Du vill förse BMP-bilderna med en RLE-kodning (Run-Length Encoding).  
Läge  
I detta område väljer Du läge för export.  
Original  
Klicka här om Du vill behålla originalläget.  
Upplösning  
Klicka här om Du vill spara bilden med en bestämd upplösning.  
I listrutan hittar Du de upplösningar som finns tillgängliga.  
Storlek  
Klicka här om Du vill spara bilden med en bestämd storlek.  
Bredd  
I detta rotationsfält ställer Du in bredden.  
Höjd  
Här definierar Du höjden.  
Mer information om filtrering finns i avsnittet om import - och exportfilter.  
GIF-alternativ  
I den här dialogrutan gör du inställningar för export av filer i GIF-format.  
Läge  
I det här området hittar du kryssrutan Interlaced.  
Interlaced  
Välj den här rutan om du vill använda sammanflätning (Interlaced=sammanflätad) vid exporten.  
Detta rekommenderas vid stora GIF-bilder eftersom du då kan se hela bilden innan laddningen är klar.  
Ritobjekt  
I det här området finns rutan Spara transparent  
Spara transparent  
Markera den här rutan om bildens bakgrund ska sparas transparent.  
I en GIF-bild syns då bara objekten.  
Du definierar den färg i bilden som ska vara transparent med hjälp av Pipett.  
Det finns mer information om filtrering i avsnittet om import - och exportfilter.  
Dif-import / export / Lotusimport / DBaseimport  
Här väljer Du ut alternativ för export resp. import.  
De här dialogerna visas automatiskt när Du väljer motsvarande filtyp.  
Teckenuppsättning  
Välj den teckenuppsättning som ska användas vid export respektive import i listrutan.  
Det finns mer information om filtrering i avsnittet Information om import - och exportfilter.  
Textexport  
I den här dialogrutan väljer du alternativ för textexporten.  
Dialogrutan visas om du använder filtypen "Text CSV" när du sparar tabelldata och har markerat rutan Redigera filterinställningar i dialogrutan Spara som.  
Fältalternativ  
I det här området bestämmer du vilken fältdelare, textavgränsare, och vilken teckenuppsättning som ska användas för textexporten.  
Teckenuppsättning  
I det här kombinationsfältet väljer du teckenuppsättning.  
Fältavgränsare  
Välj den fältavgränsare som står mellan två datafält.  
Textavgränsare  
Här väljer du textavgränsaren som omsluter alla datafält av typen text.  
Mer information om filtrering finns i avsnittet Information om import - och exportfilter.  
Textimport  
Välj här alternativen för import av data från en textfil med fältavgränsare.  
Import  
I detta område väljer Du från och med vilken rad Du vill överta data och i vilken teckenuppsättning informationen har sparats.  
Från rad  
I detta rotationsfält anger Du den första rad från vilken data ska övertas.  
Raderna visas i förhandsvisningsfönstret nederst i dialogrutan.  
I de flesta fall vill Du förmodligen inte importera den första raden om kolumnhuvudena finns där.  
Teckenuppsättning  
I det här kombinationsfältet väljer du den teckenuppsättning i vilken de data som ska importeras har sparats.  
Delningsalternativ  
I området för delningsalternativ väljer du om datafälten i textfilen ska skiljas åt med fältavgränsare eller om datafälten ska ha fasta bredder.  
Fast bredd  
Välj det här alternativet om datafälten i texten bara är åtskilda från varandra med sin bredd.  
Du ställer sedan in datafältens bredd i förhandsvisningsfönstret med musen.  
Klicka på fönstrets linjal och flytta markeringspunkten dit du vill ha den.  
Delad  
Välj det här alternativet om datafälten i texten är separerade med fältavgränsare.  
Tabulator  
Välj det här alternativet om datafälten är tabbavgränsade.  
Semikolon  
Välj det här alternativet om datafälten är separerade med semikolon.  
Komma  
Välj det här alternativet om datafälten är separerade med kommatecken.  
Blanksteg  
Välj det här alternativet om datafälten är separerade med blanksteg.  
Andra  
Välj det här alternativet om datafälten är separerade med något annat tecken.  
Skriv tecknet i det högra textfältet.  
Sammanfatta fältavgränsare  
Välj det här alternativet om flera på varandra följande fältavgränsare ska sammanfogas till en enda fältavgränsare.  
Detta påverkar direkt importen av tomma datafält.  
Textavgränsare  
I det här kombinationsfältet väljer du de avgränsningstecken som kan rama in enskilda datafält, om fältavgränsningstecknet förekommer i dem.  
Dessa textavgränsare måste vara angivna redan när textfilen skapas.  
Du kan ange tecknet direkt.  
Fält  
I ett förhandsvisningsfönster visas effekten av de inställningar Du gör.  
Typ  
I kombinationsfältet Typ väljer du i vilken typ datafältet i den kolumn som markerats i förhandsvisningsfönstret ska importeras.  
Välj bland följande alternativ:  
Typ  
Funktion  
Standard  
%PRODUCTNAME avgör själv typen.  
Text  
Tecknen övertas oförändrat som text.  
Datum (DMÅ)  
Tecken övertas som datum (Dag, Månad, År).  
Datum (MDÅ)  
Tecken övertas som datum (Månad, Dag, År).  
Datum (ÅMD)  
Tecken övertas som datum (År, Månad, Dag).  
Engelska (US)  
Något sifferformat ställs då inte in.  
Poster som inte innehåller några tal formaterade enligt amerikansk standard behandlas som under Standard.  
dölj  
Tecknen övertas inte.  
När Du importerar sifferfält som kan inledas med en eller flera nollor (telefonnummer, postnummer) ger Du dem typen Text.  
Förhandsvisning  
I området Förhandsvisning visas ett exempel på hur många tecken i en datapost som övertas i kolumnen (datafältet).  
Här kan du markera kolumner och sedan tilldela dem en typ i kombinationsfältet Typ.  
I samband med Fast bredd kan du även ställa in datafältens bredd i förhandsvisningsfönstret.  
I kombinationsfältet Typ väljer du "Dölja".  
Mer information om filter finns i Information om import - och exportfilter.  
Varning - Utskriftsalternativ  
Den här dialogrutan öppnas om sidinställningarna inte stämmer överens med det utskriftsområde som Du har definierat.  
Detta kan t ex hända om Du har ritat en rektangel som är större än det sidformat som Du har valt.  
Utskriftsalternativ  
Anpassa sidan till utskriftsområdet  
Klicka här för att anpassa sidan till utskriftsområdet.  
Utskriftsområdet styrs av det pappersformat som Du har valt.  
Om Du väljer det här alternativet visas inte dialogrutan Varning - Utskriftsalternativ när Du skriver ut i fortsättningen.  
Skriv ut på flera sidor  
Klicka här om Du vill fördela utskriften över flera sidor.  
Utskriftsområdet för t ex en alltför stor rektangel delas upp på flera sidor.  
Klipp  
Om Du väljer det här alternativet kapas allt som ligger utanför det tillgängliga utskriftsområdet bort och tas inte med i utskriften.  
PNG-alternativ  
Här väljer du kompressionsförhållande och Interlaced-läge när du sparar en bild som PNG.  
Kompression 0..9  
I detta rotationsfält väljer Du kompressionsvärde för grafiken, från 0 (ingen kompression) till 9 (maximal kompression).  
Ju högre kompressionsvärde desto mer datortid krävs, samtidigt som resultatet kräver något mindre antal byte.  
Interlaced  
Markera det här fältet om grafiken ska sparas i Interlaced-läge.  
EPS exportalternativ  
Här kan du definiera olika alternativ för exporten.  
Du kan skriva ut din fil med en Post Script-skrivare.  
Med andra skrivare skrivs förhandsvisningen ut.  
Förhandsvisning  
I det här området definierar du om du vill ha en förhandsvisning eller inte.  
Förhandsvisning bild (TIF)  
Markera detta fält om en förhandsvisningsgrafik i TIF-format ska exporteras tillsammans med den egentliga PostScript-filen.  
Interchange (EPSI)  
Markera det här fältet om ett monokromt förhandsvisningsgrafikobjekt i EPSI-format ska exporteras tillsammans med den egentliga PostScript-filen.  
Detta format innehåller bara utskrivbara tecken i 7-bitars ASCII-kod.  
Version  
I området Version bestämmer du dig för en PostScript-nivå.  
Nivå 1  
På den här nivån är inte någon komprimering tillgänglig.  
Välj det här alternativet om din PostScript-skrivare inte stöder nivå 2.  
Nivå 2  
Det här alternativfältet väljer du om din skrivare kan skriva ut såväl bitmaps i färg och palettgrafik som komprimerad grafik.  
Färgformat  
Alternativen i området Färgformat låter dig välja mellan export i färg eller i gråskalor.  
Färg  
Det här alternativfältet aktiverar du om din fil ska exporteras med färger.  
Gråskalor  
Om du väljer det här alternativet exporteras filen i gråskalor.  
Kompression  
I det här området väljer du om filen ska exporteras komprimerat.  
LZW-kodning  
LZW är förkortningen för "Lempel Ziv Welch" vilket är namnen för upphovsmännen till denna komprimeringsalgoritm.  
Om du vill använda den, aktiverar du alternativfältet.  
Ingen  
Om ingen komprimering ska användas, väljer du det här alternativet.  
Textinställningar  
Här väljer du om text exporteras med eller utan information om konturformen för varje enskilt tecken.  
Urval  
Effekt  
Exportera alltid glyfkonturer  
I förinställningen exporteras tecknens former.  
Exportera aldrig glyfkonturer  
Med den här inställningen exporteras inte formerna.  
PBM / PPM / PGM alternativ  
Välj här i vilket format filen ska exporteras.  
Den här dialogrutan visas vid export i formatet Portable Bitmap (PBM), Portable Pixelmap (PPM) och Portable Greymap (PGM).  
Filtyp  
Här väljer Du format för exporten av filen.  
Binär  
Här väljer Du export i binärformat.  
Den skapade filen är mindre än en text (ASCII )-fil.  
Text  
Här markerar Du om Du vill genomföra exporten i textformat, det vill säga ASCII -format.  
En sådan fil är större än en binär.  
ASCII filteralternativ  
Välj här med vilka alternativ (standardteckensnitt, språk, teckenuppsättning, brytning) textdokumentet ska importeras resp. exporteras.  
Dialogrutan visas så snart du laddar eller sparar en ren ascii-fil utan att ange ett annat filter.  
Filtret heter "Text - kodad".  
Egenskaper  
I området egenskaper gör du inställningar för import eller export av din fil.  
Du kan definiera vilken teckenuppsättning, vilket standardteckensnitt, vilket språk och vilken styckebrytning som ska användas.  
Vid export går det dock bara att bestämma teckenuppsättningen och styckebrytningen.  
Teckenuppsättning  
Här kan du välja bland olika teckenuppsättningar som till exempel System eller Unicode.  
Standardteckensnitt  
Med inställningen av ett standardteckensnitt definierar du om texten ska visas i t.ex. Arial eller Times New Roman.  
Det går bara att välja standardteckensnitt vid import.  
De teckensnitt som är tillgängliga på din dator visas.  
Språk  
Här kan du ställa in språket i texten om det inte redan är inställt.  
Det är bara möjligt att göra den här inställningen vid import.  
Styckebrytning  
CR står för "Carriage Return" och LF för "Linefeed ".  
De här termerna kommer från den tiden när man använde elektroniska skrivmaskiner.  
CR & LF  
Alternativet skapar både en "Carriage Return" och en "Linefeed ".  
I standardinställningen är fältet aktiverat.  
CR  
Använd det här alternativet om du vill att bara en "Carriage Return" ska skapas.  
LF  
Aktivera det här fältet om du vill att en "Linefeed" ska skapas.  
Meny Arkiv  
Meny Arkiv - Nytt  
Ikon Nytt på funktionslisten (ikonen visar den aktuella dokumenttypen)  
Nytt  
Kommando Ctrl +N  
Meny Arkiv - Nytt - Mallar och dokument  
Tangentkombinationen Skift + Kommando Ctrl +N  
Meny Arkiv - Nytt - Etiketter...  
Meny Arkiv - Nytt - Etiketter... - fliken Etiketter  
Menyn Arkiv - Nytt - Etiketter... - fliken Format  
Menyn Arkiv - Nytt - Visitkort... - fliken Format  
Menyn Arkiv - Nytt - Etiketter... - fliken TillÃ¤gg  
Menyn Arkiv - Nytt - Visitkort... - fliken TillÃ¤gg  
Menyn Arkiv - Nytt - Visitkort...  
Menyn Arkiv - Nytt - Visitkort... - fliken Medium  
Menyn Arkiv - Nytt - Visitkort... - fliken Visitkort  
Menyn Arkiv - Nytt - Visitkort... - fliken Privat  
Menyn Arkiv - Nytt - Visitkort... - fliken AffÃ¤rsmÃ¤ssig  
Menyn Arkiv - Öppna...  
Tangentkombinationen Kommando Ctrl +O  
Ikon på funktionslisten:  
Öppna fil  
Menyn Arkiv - Öppna, vald filtyp Text -kodad  
Menyn Arkiv - Spara som, vald filtyp Text - kodad  
Menyn Arkiv - AutoPilot  
Meny Arkiv - AutoPilot - Brev...  
Meny Arkiv - AutoPilot - Brev... - sida 1  
Meny Arkiv - AutoPilot - Brev / Fax... - sida 2  
Meny Arkiv - AutoPilot - Brev... - sida 3  
Meny Arkiv - AutoPilot - Brev... - sida 4  
Meny Arkiv - AutoPilot - Brev... - sida 5  
Meny Arkiv - AutoPilot - Brev / Fax... sida 6  
Meny Arkiv - AutoPilot - Brev... - sida 7  
Menyn Arkiv - AutoPilot - Brev... - sida 8 / Fax... sida 7 / PM... sida 4 / Agenda... sida 5  
Menyn Arkiv - AutoPilot - Brev... - sida 9  
Menyn Arkiv - AutoPilot - Fax...  
Menyn Arkiv - AutoPilot - Fax... - sida 1  
Menyn Arkiv - AutoPilot - Fax... - sida 3  
Menyn Arkiv - AutoPilot - Fax... - sida 4  
Menyn Arkiv - AutoPilot - Fax... - sida 5  
Menyn Arkiv - AutoPilot - Fax... - sida 8  
Menyn Arkiv - AutoPilot - PM...  
Menyn Arkiv - AutoPilot - PM... - sida 1  
Menyn Arkiv - AutoPilot - PM... - sida 2  
Menyn Arkiv - AutoPilot - PM... - sida 3  
Menyn Arkiv - AutoPilot - PM... - sida 5  
Menyn Arkiv - AutoPilot - Agenda...  
Menyn Arkiv - AutoPilot - Agenda... - sida 1  
Menyn Arkiv - AutoPilot - Agenda... - sida 2  
Menyn Arkiv - AutoPilot - Agenda... - sida 3  
Menyn Arkiv - AutoPilot - Agenda... - sida 4  
Menyn Arkiv - AutoPilot - Agenda... - sida 6  
Menyn Arkiv - AutoPilot - Presentation...  
Menyn Arkiv - AutoPilot - Presentation - sida 1  
Menyn Arkiv - AutoPilot - Presentation - sida 2  
Menyn Arkiv - AutoPilot - Presentation - sida 3  
Menyn Arkiv - AutoPilot - Presentation - sida 4  
Menyn Arkiv - AutoPilot - Presentation - sida 5  
Menyn Arkiv - AutoPilot - Web - sida...  
Menyn Arkiv - AutoPilot - FormulÃ¤r  
Menyn Arkiv - AutoPilot - FormulÃ¤r - Databasurval  
Menyn Arkiv - AutoPilot - FormulÃ¤r - Utformning  
Formulärutkast - klicka på ikonen Grupperingsram på utrullningslisten Formulärfunktioner och rita upp en ram  
Formulärutkast - klicka på ikonen Grupperingsram på utrullningslisten Formulärfunktioner och rita upp ram - AutoPilot sida 1  
Formulärutkast - klicka på ikonen Grupperingsram på utrullningslisten Formulärfunktioner och rita upp en ram - AutoPilot sida 2  
Formulärutkast - klicka på ikonen Grupperingsram på utrullningslisten Formulärfunktioner och rita upp en ram - AutoPilot sida 3  
Formulärutkast - klicka på ikonen Grupperingsram på utrullningslisten Formulärfunktioner och rita upp en ram - AutoPilot sida 4.  
Det måste redan finnas en databaskoppling.  
Formulärutkast - klicka på ikonen Grupperingsram på utrullningslisten Formulärfunktioner och rita upp en ram - sista sidan i AutoPiloten  
Menyn Arkiv - AutoPilot - Dokumentkonverterare  
Menyn Arkiv - AutoPilot - Dokumentkonverterare  
Menyn Arkiv - AutoPilot - Dokumentkonverterare  
Menyn Arkiv - AutoPilot - %PRODUCTNAME 5.2 databasimport  
Menyn Arkiv - AutoPilot - %PRODUCTNAME 5.2 databasimport - Definiera källa  
Menyn Arkiv - AutoPilot - %PRODUCTNAME 5.2 databasimport - Element som ska importeras  
Menyn Arkiv - AutoPilot - %PRODUCTNAME 5.2 databasimport - Anpassa sökväg  
Menyn Arkiv - AutoPilot - %PRODUCTNAME 5.2 databasimport - Formulärimport  
Menyn Arkiv - AutoPilot - %PRODUCTNAME 5.2 databasimport - Sökningsimport  
Menyn Arkiv - AutoPilot - %PRODUCTNAME 5.2 databasimport - Sammanfattning  
Menyn Arkiv - AutoPilot - Eurokonverterare...  
AutoPilot Adressdatakälla (startar automatiskt första gången %PRODUCTNAME startas)  
Menyn Arkiv - AutoPilot - Adressdatakälla  
AutoPilot för adressdatakällor - Ytterligare inställningar  
AutoPilot för adressdatakällor - Välj tabell  
AutoPilot för adressdatakällor - Datakällrubrik  
AutoPilot för adressdatakällor - Fälttilldelning  
Menyn Arkiv - Stäng  
Menyn Arkiv - Spara  
Tangentkombinationen Kommando Ctrl +S  
Ikon på funktions - eller databaslisten:  
Spara dokument  
Välj GIF som filtyp, dialogrutan öppnas automatiskt  
Välj PNG som filtyp, dialogrutan öppnas automatiskt  
Välj BMP som filtyp, dialogrutan öppnas automatiskt  
Välj JPEG som filtyp, dialogrutan öppnas automatiskt  
Den här dialogrutan öppnas automatiskt  
Välj Webbsida som filtyp, sidan 1 i AutoPiloten  
Välj Webbsida som filtyp, sidan 2 i AutoPiloten  
Välj Webbsida som filtyp, sidan 3 i AutoPiloten  
Välj Webbsida som filtyp, sidan 4 i AutoPiloten  
Välj Webbsida som filtyp, sidan 5 i AutoPiloten  
Välj Webbsida som filtyp, sidan 6 i AutoPiloten  
Välj SVM / WMF / PICT / MET som filtyp, dialogrutan öppnas automatiskt  
Menyn Arkiv - Spara allt  
Menyn Arkiv - Spara som...  
Menyn Arkiv - Ladda på nytt  
Menyn Arkiv - Egenskaper...  
Menyn Arkiv - Egenskaper... - fliken Allmänt  
Menyn Arkiv - Egenskaper... - fliken Beskrivning  
Menyn Arkiv - Egenskaper... - fliken Användare  
Menyn Arkiv - Egenskaper... - fliken Statistik  
Menyn Arkiv - Egenskaper... - fliken Internet  
Menyn Arkiv - Dokumentmall  
Menyn Arkiv - Dokumentmall - Förvalta  
Meny Arkiv - Dokumentmall - Administrera, kommandoknapp Adressbok  
Menyn Arkiv - Dokumentmall - Adressbokskälla  
Menyn Arkiv - Dokumentmall - Adressbokskälla, sedan kommandoknapp Administrera  
Menyn Verktyg - Datakällor Menyn Verktyg - Datakällor  
Menyn Arkiv - Dokumentmall - Spara  
Menyn Arkiv - Dokumentmall - Redigera  
Menyn Arkiv - Förhandsgranskning  
Menyn Arkiv - Skrivarinställning...  
Menyn Arkiv - Dokumentmall... - Förvalta...  
Kommandon - Skrivarinställningar...  
Menyn Arkiv - AutoPilot - Brev - sidan 9  
Menyn Arkiv - Skicka  
Menyn Arkiv - Skicka - Dokument som e-post...  
Menyn Arkiv - Dokument som e-post...  
Menyn Arkiv - Skicka - Skapa samlingsdokument  
Menyn Arkiv - Skriv ut...  
Tangentkombinationen Kommando Ctrl +P  
Ikon på funktionslisten:  
Skriv ut fil direkt  
Ikon på förhandsgranskningslisten i ett textdokument:  
Skriv ut förhandsgranskning  
Menyn Arkiv - Avsluta  
Tangentkombinationen Kommando Ctrl +Q  
Menyn Arkiv - Nytt - Samlingsdokument  
Välj filtyp: "Text CSV"  
Välj EPS som filtyp, dialogrutan öppnas automatiskt  
Menyn Arkiv - Exportera..., välj PBM, PPM eller PGM som filtyp, dialogrutan öppnas automatiskt  
Menyn Arkiv - Versioner  
Menyn Redigera  
Menyn Redigera - Ångra  
Tangentkombinationen Kommando Ctrl +Z  
Ikon på funktions - eller databaslisten:  
Ångra  
Menyn Redigera - Återställ  
Ikon på funktionslisten:  
Återställ  
Menyn Redigera - Senaste kommando  
Menyn Redigera - Klipp ut  
Tangentkombinationen Kommando Ctrl +X  
Ikon på funktionslisten:  
Klipp ut  
Menyn Redigera - Kopiera  
Tangentkombinationen Kommando Ctrl +C  
Ikon på funktionslisten:  
Kopiera  
Menyn Redigera - Klistra in  
Tangentkombinationen Kommando Ctrl +V  
Ikon på funktionslisten:  
Klistra in  
Menyn Redigera - Klistra in innehÃ¥ll...  
Menyn Redigera - Markera allt  
Tangentkombinationen Kommando Ctrl +A  
Markera allt  
Menyn Redigera - Ã„ndringar  
Menyn Redigera - Ã„ndringar - Registrera  
Menyn Redigera - Ändringar - Visa Menyn Redigera - Ã„ndringar - Visa...  
Menyn Redigera - Ã„ndringar - Acceptera eller ignorera...  
Menyn Redigera - Ändringar - Acceptera eller ignorera... fliken Lista  
Menyn Format - AutoFormat - Använd och redigera ändringar - dialog AutoFormat - kommandoknapp Redigera ändringar - fliken Lista  
Menyn Redigera - Ändringar - Acceptera eller ignorera... fliken Filter  
Menyn Redigera - Ã„ndringar - Sammanfoga dokument...  
Menyn Redigera - JÃ¤mfÃ¶r dokument...  
Menyn Redigera - Ändringar - Kommentar...  
Ändra kommentar  
Menyn Redigera - Sök och ersätt...  
Tangentkombinationen Kommando Ctrl +G  
Ikon på verktygslisten (text-, tabelldokument):  
Sökning på / av  
Menyn Redigera - Sök och ersätt... - kommandoknapp Attribut...  
Menyn Redigera - Sök och ersätt... - kommandoknapp Format...  
Menyn Redigera - Sök och ersätt... - fältet Likhetssökning markerat och kommandoknappen... vald  
Vy i en databastabell: ikon Genomsök... på databaslisten - fältet Likhetssökning markerat och kommandoknappen... vald  
Formulärvy: ikon Datapostsökning på formulärlisten - fältet Likhetssökning markerat och kommandoknappen... vald  
Menyn Redigera - Navigator  
Tangent F5  
Ikon på funktionslisten:  
Navigator på / av  
Menyn Verktyg - Litteraturdatabas  
Menyn Redigera - LÃ¤nkar...  
Menyn Redigera - Länkar - Ändra länk (bara för DDE-länk)  
Markera en ram, välj sedan Redigera - Objekt - Egenskaper... - Ram - fliken Egenskaper  
Snabbmeny till en markerad ram, menykommando Egenskaper  
Menyn Redigera - PlugIn  
Menyn Redigera - Image map samt i snabbmenyn för ett markerat objekt  
Menyn Redigera - Image map, markera sedan ett område Egenskaper - Beskrivning  
Menyn Redigera - Objekt  
Menyn Redigera - Objekt - Redigera och i snabbmenyn till ett markerat objekt  
Menyn Redigera - Objekt - Ã–ppna  
Menyn Visa  
Menyn Visa - Skala...  
Zooma även med +, -, × och ÷ på det numeriska tangentbordet Zooma Ã¤ven med +, -, Ã— och Ã· pÃ¥ det numeriska tangentbordet  
Dubbelklicka på fältet 100% på statuslisten  
Meny Visa - Symbollister - Redigera  
Snabbmeny Redigera  
Meny Visa - Symbollister - Funktionslist  
Meny Visa - Symbollister - Objektlist  
Meny Visa - Symbollister - Verktygslist  
Meny Visa - Statuslist  
Menyn Visa - Symbollister - FÃ¤rglist  
Hyperlänklist - ikon Hyperlänkdialog - Internet  
Hyperlänklist - ikon Hyperlänk-dialog - fliken E-post & nyheter  
Hyperlänklist - ikon Hyperlänkdialog - Dokument  
Hyperlänklist - ikon Hyperlänkdialog - Nytt dokument  
Menyn Visa - Hela bildskärmen  
Tangent Skift + Kommando Ctrl +J  
Om ett text - eller tabelldokument är öppet:  
Menyn Visa - Datakällor  
Tangent F4  
Datakällor  
Menyn Visa - HTML-källtext  
Snabbmeny i HTML-dokument  
Visa HTML-källtext  
Meny Infoga  
Meny Infoga - Anteckning  
Meny Infoga - Skanna  
Meny Infoga - Skanna - Välj källa... (teckningsdokument, (textdokument)  
Meny Arkiv - Skanna - Välj källa... (bilddokument)  
Meny Infoga - Skanna - Rekvirera... (teckningsdokument), (textdokument)  
Meny Arkiv - Skanna - Rekvirera... (bilddokument)  
Meny Infoga - Specialtecken...  
Meny Format - Numrering / punktuppställning... - Alternativ, kommandoknapp Tecken  
Menyn Format - Numrering / punktuppställning... - Alternativ, kommandoknappen Tecken  
Ikon på utrullningslisten Infoga på verktygslisten (inte för diagram):  
Infoga specialtecken  
Meny Infoga - Objekt  
Meny Infoga - Objekt - OLE-objekt...  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga OLE-objekt  
Meny Infoga - Objekt - Plug-in...  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga plug-in  
Menyn Infoga - Objekt - Ljud...  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga ljud-plug-in  
Menyn Infoga - Objekt - Video....  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga video-plug-in  
Menyn Infoga - Objekt - Applet...  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga applet  
Menyn Infoga - Objekt - Formel...  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga %PRODUCTNAME Math-objekt Infoga Formel  
Menyn Format - AutoFormat... - AutoFormat Diagram - sida 1 av 3  
Menyn Infoga - Objekt - Diagram - AutoFormat Diagram - sida 2 av 4  
Menyn Format - AutoFormat... - AutoFormat Diagram - sida 2 av 3  
Menyn Infoga - Objekt - Diagram - AutoFormat Diagram - sida 3 av 4  
Menyn Format - AutoFormat... - AutoFormat Diagram - sida 3 av 3  
Menyn Infoga - Objekt - Diagram - AutoFormat Diagram - sida 4 av 4  
Menyn Infoga - Objekt - Diagram  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga diagram  
Menyn Infoga - Grafik - Från fil...  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga grafik  
Menyn Arkiv - Nytt - Bild  
Menyn Infoga - Ram  
Ikon på utrullningslisten Infoga objekt på verktygslisten:  
Infoga ramteknik  
Menyn Infoga - Ramteknik, efter val av en fil  
Meny - Visa - Symbollister - Hyperlänklist  
Ikon på verktygslisten (text-, tabelldokument):  
Hyperlänklist på / av  
Meny Verktyg  
Meny Verktyg - Gallery eller ikon på funktionslisten:  
Gallery  
Meny Verktyg - Gallery eller ikon på funktionslisten - kommandoknapp Nytt tema - fliken Filer  
Dialogrutan visas bara om rättstavningskontrollen hittar ett fel:  
Meny Verktyg - Rättstavning - Kontrollera...  
Tangenten F7  
Ikon på verktygslisten:  
Rättstavning  
Meny Verktyg - RÃ¤ttstavning  
Meny Verktyg - Rättstavning - Kontrollera - (dialogrutan visas bara om rättstavningskontrollen hittar ett fel) och sedan klickar du på Alternativ  
Meny Verktyg - Synonymordlista...  
Meny Verktyg - Rättstavning - Kontrollera - Synonymordlista  
Kortkommandot Kommando Ctrl +F7  
Meny Verktyg - Pipett (%PRODUCTNAME Draw und %PRODUCTNAME Impress)  
Meny Verktyg - Makro  
Meny Verktyg - Makro - Administrera - fliken Bibliotek - LÃ¶senord  
Meny Verktyg - Anpassa  
Menyn Verktyg - Anpassa - fliken Meny  
Meny Verktyg - Anpassa - fliken Tangentbord  
Menyn Verktyg - Anpassa - fliken Statuslist  
Menyn Verktyg - Anpassa... - fliken Symbollister  
Menyn Verktyg - Anpassa... - fliken Symbollister - Redigera...  
Visa - Symbollister - Redigera...  
Snabbmenyn för symbollister Redigera...  
Menyn Verktyg - Anpassa - fliken HÃ¤ndelser  
Menyn Verktyg - AutoKorrigering / AutoFormat  
Menyn Verktyg - AutoKorrigering / AutoFormat - fliken Alternativ  
Menyn Verktyg - AutoKorrigering / AutoFormat - fliken ErsÃ¤ttning  
Menyn Verktyg - AutoKorrigering / AutoFormat - fliken Undantag  
Menyn Verktyg - AutoKorrigering / AutoFormat - fliken Typografiska anfÃ¶ringstecken  
Meny Verktyg - AutoKorrigering / AutoFormat - fliken Ordkomplettering  
Menyn Verktyg - Alternativ - Tabelldokument - Vy  
Menyn Verktyg - Alternativ - Presentation / Teckning - Vy  
Menyn Verktyg - Alternativ - Teckning - AllmÃ¤nt  
Kommandoknapp för val av sökväg i diverse AutoPiloter  
Redigera -kommandoknapp för en del poster i Verktyg - Alternativ - %PRODUCTNAME - SÃ¶kvÃ¤gar  
Menyn Verktyg - Alternativ  
Menyn Verktyg - Alternativ - %PRODUCTNAME  
Menyn Verktyg - Alternativ - %PRODUCTNAME - AnvÃ¤ndardata  
Menyn Verktyg - Alternativ - %PRODUCTNAME - AllmÃ¤nt  
Menyn Verktyg - Alternativ - %PRODUCTNAME - Arbetsminne  
Menyn Verktyg - Alternativ - %PRODUCTNAME - Vy  
Menyn Verktyg - Alternativ - %PRODUCTNAME - HjÃ¤lpprogram  
Menyn Verktyg - Alternativ - %PRODUCTNAME - Skriv ut  
Menyn Verktyg - Alternativ - %PRODUCTNAME - Sökvägar  
Menyn Redigera - AutoText - Sökväg...  
Menyn Verktyg - Alternativ - %PRODUCTNAME - Färger  
Menyn Format - Yta... - fliken FÃ¤rger  
Menyn Verktyg - Alternativ - %PRODUCTNAME - Färger - Redigera  
Menyn Format - Yta... - fliken FÃ¤rger - Redigera...  
Menyn Format - 3D-effekter - ikon på fliken Belysning:  
Välj färg i färgdialogruta  
Menyn Verktyg - Alternativ - %PRODUCTNAME - TeckensnittsersÃ¤ttning  
Menyn Verktyg - Alternativ - %PRODUCTNAME - SÃ¤kerhet  
Menyn Verktyg - Alternativ - Ladda / spara  
Menyn Verktyg - Alternativ - Allmänt - sidan Spara  
Menyn Verktyg - Alternativ - Ladda / spara - VBA-egenskaper  
Menyn Verktyg - Alternativ - Ladda / Spara - Microsoft Office  
Menyn Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet  
Menyn Verktyg - Alternativ - SprÃ¥kinstÃ¤llningar  
Menyn Verktyg - Alternativ - SprÃ¥kinstÃ¤llningar - SprÃ¥k  
Menyn Verktyg - Alternativ... - Allmänt - sidan Lingvistik  
Menyn Verktyg - Alternativ - Språkinställningar - Lingvistik, välj en språkmodul i listrutan Tillgängliga språkmoduler, sedan kommandoknapp Redigera  
Menyn Verktyg - Alternativ - Språkinställningar - SÃ¶kalternativ fÃ¶r japanska  
Menyn Verktyg - Alternativ - Språkinställningar - Asiatisk layout  
Menyn Verktyg - Alternativ - Internet  
Menyn Verktyg - Alternativ... - Internet - sidan Proxy  
Menyn Verktyg - Alternativ - Internet - sidan SÃ¶kning  
Menyn Verktyg - Alternativ - Textdokument  
Menyn Verktyg - Alternativ - Textdokument - AllmÃ¤nt  
Menyn Verktyg - Alternativ - Textdokument - AllmÃ¤nt - Objekturval - kommandoknapp...  
Menyn Verktyg - Alternativ - Textdokument / HTML-dokument - Vy  
Menyn Verktyg - Alternativ - Textdokument / HTML-dokument - FormateringshjÃ¤lp  
Menyn Verktyg - Alternativ - Text - / Tabelldokument / HTML-dokument - Raster  
Menyn Verktyg - Alternativ - Textdokument - Standardteckensnitt  
Menyn Verktyg - Alternativ - Textdokument / HTML-dokument / Tabelldokument - Skriv ut  
Menyn Verktyg - Alternativ - Textdokument / HTML-dokument - Tabell  
Menyn Verktyg - Alternativ - Textdokument - Ã„ndringar  
Meny Verktyg - Alternativ - HTML-dokument  
Menyn Verktyg - Alternativ - HTML-dokument - KÃ¤lltext  
Menyn Verktyg - Alternativ - HTML-dokument - Bakgrund  
Menyn Verktyg - Alternativ - Tabelldokument  
Menyn Verktyg - Alternativ - Tabelldokument - AllmÃ¤nt  
Menyn Verktyg - Alternativ - Tabelldokument - Vy  
Menyn Verktyg - Alternativ - Tabelldokument - BerÃ¤kna  
Menyn Verktyg - Alternativ - Tabelldokument - Sorteringslistor  
Menyn Verktyg - Alternativ - Tabelldokument - Sorteringslistor - Kopiera  
Menyn Verktyg - Alternativ - Tabelldokument - Ã„ndringar  
Menyn Verktyg - Alternativ - Presentation  
Menyn Verktyg - Alternativ - Presentation / Teckning - AllmÃ¤nt  
Menyn Verktyg - Alternativ - Presentation / Teckning - Vy  
Menyn Verktyg - Alternativ - Presentation / Teckning - Raster  
Menyn Verktyg - Alternativ - Presentation / Teckning - Skriv ut  
Menyn Verktyg - Alternativ - Teckning  
Menyn Verktyg - Alternativ - Formel  
Menyn Verktyg - Alternativ - Formel - InstÃ¤llningar  
Menyn Verktyg - Alternativ - Diagram  
Menyn Verktyg - Alternativ - Diagram - GrundfÃ¤rger  
Menyn Verktyg - Alternativ - DatakÃ¤llor  
Menyn Verktyg - Alternativ - DatakÃ¤llor - FÃ¶rbindelser  
Menyn Fönster  
Menyn FÃ¶nster - Nytt fÃ¶nster  
Menyn Fönster - Förteckning över öppnade dokument  
Menyn Hjälp  
Menyn HjÃ¤lp - InnehÃ¥ll  
Menyn Hjälp - Om %PRODUCTNAME...  
Automatiskt andra gången %PRODUCTNAME startas  
Menyn Hjälp - Registrering (direkt till webbsidan)  
Symbollister  
Menyn Data - Filter - Standardfilter...  
Visning av en databastabell: ikonen Standardfilter på databaslisten  
Formulärvy: ikonen Standardfilter på formulärlisten  
Standardfilter  
Databas  
Verktyg - Datakällor - fliken Tabeller  
Verktyg - Datakällor - fliken SÃ¶kningar  
Verktyg - Datakällor - fliken LÃ¤nkar  
Meny Arkiv - Dokumentmall - Adressbokskälla, sedan kommandoknappen Administrera, sedan fliken AllmÃ¤nt  
Verktyg - Datakällor - fliken ODBC, eller så valdes databastypen Adressbok  
Kommandoknapp för val av sökväg i diverse AutoPiloter / Redigera kommandoknapp för några poster under Verktyg - Alternativ - %PRODUCTNAME - SÃ¶kvÃ¤gar  
Verktyg - Datakällor - fliken ODBC  
Välj Verktyg - Datakällor - Allmänt - databastyp Adressbok, välj LDAP adressbok så visas fliken LDAP  
Verktyg - Datakällor - fliken JDBC  
Verktyg - Datakällor - fliken dBase  
Verktyg - Datakällor - fliken dBase - Index  
Verktyg - Datakällor - fliken Text  
Verktyg - Datakällor - fliken Adabas D  
Verktyg - Datakällor - fliken ADO  
Öppna databas - snabbmeny - SQL  
Öppna databas - snabbmeny till en sökningscontainer  
Öppna databas - snabbmenyn till en tabellcontainer  
Öppna databas - snabbmenyn till en tabellcontainer eller en tabell - Nytt tabellutkast eller Redigera tabell  
Öppna databas - snabbmenyn till en tabellcontainer eller en tabell - Nytt tabellutkast eller Redigera tabell - sedan Verktyg - Indexutkast eller ikon Indexutkast  
Öppna databas - snabbmeny till en sökningscontainer - Nytt sÃ¶kningsutkast  
Öppna databas - snabbmeny till en sökningscontainer - Nytt sökningsutkast / Öppna databas - öppna sökningscontainer - snabbmeny till en sökning - Redigera sÃ¶kning  
Öppna databas - öppna sökningscontainer - snabbmeny till en sökning - Redigera sökning om tabeller eller fält i sökningen inte längre existerar.  
Öppna sökningsutkast och dubbelklicka på en förbindelselinje som ligger mellan två tabeller  
Öppna databas - snabbmenyn till en sökningscontainer eller en sökning - Nytt - Sökning - Sökningsutkast Öppna databas - snabbmenyn till en tabellcontainer eller en tabell - Nytt - Tabellvy (inte vid dBase-databaser) ikon på sökningslisten i sökningsutkastet och - vid relationsdatabassystem - i relationsfönstret:  
Lägg till tabell...  
Klicka på ikonen i relationsfönstret om det innehåller minst 2 tabeller:  
Ny relation...  
Ikon Sök datapost på databaslisten och formulärlisten  
Sök datapost...  
Ikon Sortera på databaslisten och formulärlisten  
Sortera...  
Verktyg - Datakällor - fliken Allmänt  
Datakällvy: dra-och-släpp av en sökning eller tabell till en söknings - eller tabellcontainer  
Öppna databas - snabbmeny till en formulärcontainer eller ett formulär - Nytt - Formulär  
Öppna databas - snabbmeny till en tabellcontainer - Användarinställningar  
Öppna databas - snabbmeny till en tabellcontainer - Relationer  
Urval av "Adabas D"  
Menyn Format  
Menyn Format - Standard  
Menyn Format - Tecken  
Ikon på objektlisten med textmarkören i ett objekt:  
Teckenattribut  
Menyn Format - Tecken... - fliken Teckensnitt  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Teckensnitt  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Teckensnitt  
Menyn Redigera - Sök och ersätt... - Format... - fliken Teckensnitt  
Radhuvudets snabbmeny i en öppnad databastabell - Tabellformatering... - fliken Teckensnitt  
Menyn Format - Cell... - fliken Teckensnitt (tabelldokument)  
Menyn Format - Titel - fliken Tecken (diagramdokument)  
Menyn Format - Förklaring... - fliken Tecken (diagramdokument)  
Menyn Format - Axel - fliken Tecken (diagramdokument)  
Menyn Format - Sida - Sidhuvud / Sidfot - kommandoknapp Redigera (tabelldokument)  
Snabbmenyn Teckensnitt  
Menyn Format - Tecken... - fliken Teckeneffekt  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Teckeneffekter  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Teckeneffekter  
Menyn Redigera - Sök och ersätt... - Format... - fliken Teckeneffekt  
Menyn Format - Tecken - fliken Teckeneffekt (presentations-och teckningsdokument)  
Menyn Format - Sida - Sidhuvud / Sidfot - kommandoknapp Redigera (tabelldokument)  
Meny Format - Tecken - fliken Position  
Meny Format - Mallar - Katalog - Ändra / Nytt - fliken Position  
Meny Format - Stylist - snabbmeny Ändra / Nytt - fliken Position  
Meny Redigera - Sök och ersätt - Format - fliken Position  
Meny Format - Tecken - fliken Position (presentations - och teckningsdokument)  
Menyn Format - Sida - Sidhuvud / Sidfot - kommandoknapp Redigera (tabelldokument)  
Menü Format - Tecken - fliken Asiatisk layout  
Meny Format - Mallar - Katalog - Ändra / Nytt - fliken Asiatisk layout  
Meny Format - Stylist - snabbmeny Ändra / Nytt - fliken Asiatisk layout  
Meny Redigera - Sök och ersätt - Format - fliken Asiatisk layout  
Meny Format - Stycke - fliken Asiatisk typografi (inte i HTML)  
Meny Format - Cell - fliken Asiatisk typografi  
Meny Format - Mallar - Katalog - Ändra / Nytt - fliken Asiatisk typografi  
Meny Format - Stylist - snabbmeny Ändra / Nytt - fliken Asiatisk typografi  
Menyn Format - Tecken... - fliken HyperlÃ¤nk  
Menyn Infoga - Kuvert... - fliken Format - kommandoknappen Redigera - Tecken... - fliken HyperlÃ¤nk  
Menyn Infoga - Hyperlänk...  
Menyn Format - Stycke  
Ikon på objektlisten med textmarkören i ett objekt:  
Format: stycke  
Menyn Format - Stycke... - fliken Justering  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Justering  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Justering  
Menyn Redigera - Sök och ersätt... - Format... - fliken Justering  
Snabbmenyn Justering  
Menyn Format - Stycke... - fliken Indrag och avstÃ¥nd  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Indrag och avstÃ¥nd  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Indrag och avstÃ¥nd  
Menyn Redigera - Sök och ersätt... - Format... - fliken Indrag och avstÃ¥nd  
Menyn Format - Mallar - Katalog - Ändra / Nytt... - fliken Indrag och avstÃ¥nd  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Indrag och avstÃ¥nd  
Menyn Format - Stycke... - fliken Tabulator  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Tabulator  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Tabulator  
Menyn Format - Stycke... - fliken Tabulator (presentations - och tabelldokument)  
Dubbelklicka på linjallisten  
Menyn Format - Stycke... - fliken Inramning  
Menyn Format - Grafik... - fliken Inramning  
Menyn Format - Objekt... - fliken Inramning  
Menyn Format - Tabell... - fliken Inramning  
Menyn Format - Ram... - fliken Inramning  
Menyn Format - Sida... - fliken Inramning  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Inramning  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Inramning  
Menyn Format - Sida... - fliken Sidhuvud - TillÃ¤gg  
Menyn Format - Sida... - fliken Sidfot - TillÃ¤gg  
Menyn Format - Cell... - fliken Inramning  
Meny Format - Stycke - fliken Inramning AvstÃ¥nd till innehÃ¥ll  
Menyn Format - Sida - Inramning - AvstÃ¥nd till innehÃ¥ll  
Menyn Format - Stycke... - fliken Bakgrund  
Menyn Format - Tecken... - fliken Bakgrund  
Menyn Format - Grafik... - fliken Bakgrund  
Menyn Format - Tabell... - fliken Bakgrund  
Menyn Format - Ram... - fliken Bakgrund  
Menyn Format - Sida... - fliken Bakgrund  
Menyn Format - Sida... - fliken Sidhuvud - TillÃ¤gg  
Menyn Format - Sida... - fliken Sidfot - TillÃ¤gg  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Bakgrund  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Bakgrund  
Menyn Infoga eller Redigera - Område... - fliken Bakgrund  
Menyn Infoga - Kuvert... - fliken Format - kommandoknappen Redigera - Tecken... - fliken Bakgrund  
Menyn Verktyg - Alternativ... - HTML-dokument... fliken Bakgrund  
Menyn Format - Cell... - fliken Bakgrund  
Menyn Format - Sida... - fliken Administrera  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Administrera  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Administrera  
Menyn Format - Sida... - fliken Sida  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Sida  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Sida  
Menyn Format - Sida... - fliken Sidhuvud  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Sidhuvud  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Sidhuvud  
Menyn Format - Sida... - fliken Sidfot  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Sidfot  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Sidfot  
Menyn Format - Stylist  
Tangent F11  
Ikon på funktionslisten:  
Stylist  
Menyn Format - Mallar  
Menyn Format - Mallar - Katalog...  
Tangenterna Kommando Ctrl +Y  
Menyn Format - 3D-effekter  
Ikon på verktygslisten:  
Menyn Format - Mallar - Katalog...  
Menyn Format - 3D-effekter - fliken Favoriter  
Menyn Format - 3D-effekter - fliken Geometri  
Menyn Format - 3D-effekter - fliken Visning  
Menyn Format - 3D-effekter - fliken Belysning  
Menyn Format - 3D-effekter - fliken Texturer  
Menyn Format - 3D-effekter - fliken Material  
Menyn Format - Numrering / punktuppställning...  
Ikon på objektlisten:  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Justering  
Punktuppställningstecken  
Menyn Format - Numrering / punktuppställning... - fliken Alternativ  
Stylist - Presentationsobjektmallar - en dispositionsformatmalls snabbmeny Nytt... / Ã„ndra...  
Stylist - Numreringsformatmallar - snabbmenyn Nytt... / Ã„ndra...  
Menyn Format - Numrering / punktuppställning... - fliken Punkter  
Stylist - Presentationsobjektmallar - en dispositionsformatmalls snabbmeny Nytt... / Ã„ndra...  
Stylist - Numreringsformatmallar - snabbmenyn Nytt... / Ã„ndra...  
Menyn Format - Numrering / punktuppställning... - fliken Numreringstyp  
Stylist - Presentationsobjektmallar - en dispositionsformatmalls snabbmeny Nytt... / Ã„ndra...  
Stylist - Numreringsformatmallar - snabbmenyn Nytt... / Ã„ndra...  
Menyn Format - Numrering / punktuppställning... - fliken Disposition  
Stylist - Numreringsformatmallar - snabbmenyn Nytt... / Ã„ndra...  
Menyn Format - Numrering / punktuppställning... - fliken Grafik  
Stylist - Presentationsobjektmallar - en dispositionsformatmalls snabbmeny Nytt... / Ã„ndra...  
Stylist - Numreringsformatmallar - snabbmenyn Nytt... / Ã„ndra...  
Menyn Format - Numrering / punktuppställning... - fliken Position  
Menyn Verktyg - Kapitelnumrering... - fliken Position  
Stylist - Numreringsformatmallar - snabbmenyn Nytt... / Ã„ndra...  
Menyn Format - Grafik - fliken BeskÃ¤ra  
Ikon på grafikobjektlisten:  
Menyn Format - Bokstäver / tecken  
Snabbmeny (text) Bokstäver / tecken  
Menyn Format - Ruby  
Meny Format  
Klicka på ikonen Tabellkontrollfält på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Klicka på ikonen Tabellkontrollfält på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Det får inte finnas någon databasanslutning i det aktuella formuläret.  
Klicka på ikonen Tabellkontrollfält på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Det måste redan finnas en databasanslutning.  
Klicka på ikonen Kombinationsfält eller Listruta på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Det måste redan finnas en databasanslutning i det aktuella formuläret.  
Klicka på ikonen Kombinationsfält eller Listruta på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Det måste redan finnas en databasanslutning i det aktuella formuläret.  
AutoPilot - sida 1.  
Klicka på ikonen Kombinationsfält eller Listruta på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Det måste redan finnas en databasanslutning i det aktuella formuläret.  
AutoPilot - sida 2.  
Klicka på ikonen Listruta på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Det måste redan finnas en databasanslutning i det aktuella formuläret.  
AutoPilot - sida 3.  
Klicka på ikonen Kombinationsfält på utrullningslisten Formulärfunktioner på verktygslisten och rita upp ett fält med musen.  
Det måste redan finnas en databasanslutning i det aktuella formuläret.  
AutoPilot - sida 3.  
Ikon på utrullningslisten Kontrollfält i makrolisten:  
Egenskaper  
Meny Format - Formulär  
Snabbmenyn i ett markerat formulärelement Formulär...  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge:  
Formuläregenskaper  
Meny Format - Formulär - Allmänt  
Snabbmenyn i ett markerat formulärelement Formulär... - fliken Allmänt  
Ikonen Formuläregenskaper på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge - fliken Allmänt  
Meny Format - Formulär... - fliken Data  
Snabbmenyn i ett markerat formulärelement Formulär... - fliken Data  
Ikonen Formuläregenskaper på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge - fliken Data  
Menyn Format - Formulär... - fliken Händelser  
Snabbmenyn i ett markerat formulärelement Formulär... - fliken Händelser  
Ikonen Formuläregenskaper på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge - fliken Händelser  
Menyn Format - Kontrollfält  
Snabbmenyn i ett markerat formulärelement Kontrollfält...  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge:  
Kontrollfältegenskaper  
Menyn Format - Kontrollfält - fliken Allmänt  
Snabbmenyn i ett markerat formulärelement Kontrollfält... - Sida Flik Allmänt  
Ikonen Kontrollfältegenskaper på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge - fliken Allmänt  
Menyn Format - Kontrollfält... - fliken Data  
Snabbmenyn i ett markerat formulärelement Kontrollfält... - fliken Data  
Ikonen Kontrollfältegenskaper på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge - fliken Data  
Menyn Format - Kontrollfält... - fliken Händelser  
Snabbmenyn i ett markerat formulärelement Kontrollfält... - fliken Händelser  
Ikonen Kontrollfältegenskaper på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge - fliken Händelser  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge:  
Aktiveringsordningsföljd  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge:  
Lägg till fält  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge:  
Formulär Navigator  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten och på objektlisten i utkastläge:  
Utkastläge på / av  
Öppna Formulär-Navigator - Markera formulär - öppna snabbmenyn - Öppna i utkastläge  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten:  
Öppna i utkastläget  
Ikon på utrullningslisten Formulärfunktioner på verktygslisten:  
Autopilot på / av  
Menyn Format - Placering (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Snabbmeny Placering (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Meny Ändra - Placering (%PRODUCTNAME Draw)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc) eller verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Placering  
Meny Format - Placering - Längst fram (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Placering - Längst fram (%PRODUCTNAME Draw)  
Skift + Kommando Ctrl +" + "(%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Snabbmeny Placering - Längst fram (%PRODUCTNAME Impress)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc) eller verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Längst fram  
Meny Format - Placering - Längre fram (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Placering - Längre fram (%PRODUCTNAME Draw)  
Kommando Ctrl +" + "(%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Snabbmeny Placering - Längre fram (%PRODUCTNAME Impress)  
Längre fram  
Meny Format - Placering - Längre bak (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Placering - Längre bak (%PRODUCTNAME Draw)  
Kommando Ctrl +" - "(%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Snabbmeny Placering - Längre bak (%PRODUCTNAME Impress)  
Längre bak  
Meny Format - Placering - Längst bak (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Placering - Längst bak (%PRODUCTNAME Draw)  
Skift + Kommando Ctrl +" - "(%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Snabbmeny Placering - Längst bak (%PRODUCTNAME Impress)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc) eller verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Längst bak  
Meny Format - Placera - I förgrunden  
Ikon på objektlisten:  
I förgrunden  
Meny Format - Placera - I bakgrunden  
Ikon på objektlisten:  
I bakgrunden  
Meny Format - Justering (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Justering (markerade objekt) (%PRODUCTNAME Draw)  
Snabbmeny Justering (markerade objekt) (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Meny Format - Justering - Vänster (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Justering - Vänster (markerade objekt) (%PRODUCTNAME Draw)  
Snabbmeny Justering - Vänster (markerade objekt) (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc), ikon på verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Vänster (vid ram)  
Vänster (vid ritobjekt)  
Meny Format - Justering - Centrerad (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Justering - Centrerad (markerade objekt) (%PRODUCTNAME Draw)  
Snabbmeny Justering - Centrerat (markerade objekt) (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc), ikon på verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Centrerad (vid ram)  
Centrerad (vid ritobjekt)  
Meny Format - Justering - Höger  
Meny Ändra - Justering - Höger (markerade objekt) (%PRODUCTNAME Draw)  
Snabbmeny Justering - Höger (markerade objekt) (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc), ikon på verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Höger (vid ram)  
Höger (vid ritobjekt)  
Meny Format - Justering - Överst (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Justering - Överst (markerade objekt) (%PRODUCTNAME Draw)  
Snabbmeny Justering - Överst (markerade objekt) (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc), ikon på verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Överst (vid ram)  
Överst (vid ritobjekt)  
Meny Format - Justering - Mitt (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Justering - Mitt (markerade objekt) (%PRODUCTNAME Draw)  
Snabbmeny Justering - Mitten (markerade objekt) (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc), ikon på verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Vertikalt centrerad (vid ram)  
Centrerad (vid ritobjekt)  
Meny Format - Justering - Underst (%PRODUCTNAME Writer, %PRODUCTNAME Calc)  
Meny Ändra - Justering - Underst (markerade objekt) (%PRODUCTNAME Draw)  
Snabbmeny Justering - Underst (markerade objekt) (%PRODUCTNAME Impress, %PRODUCTNAME Draw)  
Ikon på objektlisten (%PRODUCTNAME Writer, %PRODUCTNAME Calc), ikon på verktygslisten (%PRODUCTNAME Impress, %PRODUCTNAME Draw):  
Vid underkant (vid ram)  
Underst (vid ritobjekt)  
Meny Format - Förankring  
Ikon på objektlisten:  
Byt förankring  
Byt förankring  
Meny Format - Förankring - Vid sidan  
Meny Format - Förankring - Vid stycke  
Meny Format - Förankring - Vid tecken  
Meny Format - Förankring - Som tecken  
Meny Format - Förankring - Till ramen  
Meny Format - Förankring - Vid cellen  
Menyn Format  
Menyn Format - Linje...  
Ikon på objektlisten:  
Linje  
Menyn Format - Linje... - fliken Linje  
Menyn Format - Formatmallar - Katalog... - Ändra / Nytt... - fliken Linje (presentationsdokument)  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Linje (presentationsdokument)  
Menyn Format - Titel - fliken Inramning (diagramdokument)  
Menyn Format - Förklaring... - fliken Inramning (diagramdokument)  
Menyn Format - Axel - fliken Linje (diagramdokument)  
Menyn Format - Gitter... - fliken Linje (diagramdokument)  
Menyn Format - Diagramvägg... - fliken Inramning (diagramdokument)  
Menyn Format - Diagramgolv... - fliken Inramning (diagramdokument)  
Menyn Format - Diagramområde... - fliken Inramning (diagramdokument)  
Menyn Format - Linje... - fliken Linjestilar  
Menyn Format - Linje... - fliken Linjeslut  
Menyn Format - Yta  
Ikon på objektlisten:  
Yta  
Menyn Format - Yta... - fliken Yta  
Menyn Format - Formatmallar - Katalog... - Ändra / Nytt... - fliken Yta (presentationsdokument)  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Yta (presentationsdokument)  
Menyn Format - Titel - fliken Yta (diagramdokument)  
Menyn Format - Förklaring... - fliken Yta (diagramdokument)  
Menyn Format - Diagramvägg... - fliken Yta (diagramdokument)  
Menyn Format - Diagramgolv... - fliken Yta (diagramdokument)  
Menyn Format - Diagramområde... - fliken Yta (diagramdokument)  
Menyn Format - Sida... - fliken Bakgrund (i %PRODUCTNAME Impress och %PRODUCTNAME Draw)  
Menyn Format - Yta... - fliken FÃ¤rger  
Menyn Verktyg - Alternativ - %PRODUCTNAME - Färger  
Menyn Format - Yta... - fliken Transparens (ritdokument)  
Menyn Format - Yta... - fliken Transparens (presentationsdokument)  
Menyn Format - Diagramvägg... - fliken Transparens (diagramdokument)  
Menyn Format - Diagramområde... - fliken Transparens (diagramdokument)  
Menyn Format - Diagramgolv... - fliken Transparens (diagramdokument)  
Menyn Format - Titel - Alla titlar.. - fliken Transparens (diagramdokument)  
Menyn Format - Titel - Huvudrubrik... - fliken Transparens (diagramdokument)  
Menyn Format - Titel - Underrubrik... - fliken Transparens (diagramdokument)  
Menyn Format - Titel - X-axeltitel... - fliken Transparens (diagramdokument)  
Menyn Format - Titel - Y-axeltitel... - fliken Transparens (diagramdokument)  
Menyn Format - Titel - X-axeltitel... - fliken Transparens (diagramdokument)  
Menyn Format - Objektegenskaper... - Datapunkt - fliken Transparens (diagramdokument)  
Menyn Format - Objektegenskaper... - Dataserie - fliken Transparens (diagramdokument)  
Menyn Format - Yta... - fliken Skugga  
Menyn Format - Yta... - fliken FÃ¤rggradienter  
Menyn Format - Yta... - fliken Skrafferingar  
Menyn Format - Yta... - fliken BitmapmÃ¶nster  
Menyn Format - Text  
Meny Format - Text... - fliken Text  
Meny Format - Text... - fliken Animerad text  
Menyn Format - Position och storlek...  
F4 F4  
Ikon på objektlisten vid markerat kontrollfält:  
Position och storlek  
Menyn Format - Position och storlek... - fliken Position  
Menyn Format - Position och storlek... - fliken Storlek  
Menyn Format - Position och storlek... - fliken Rotation  
Ikon på objektlisten:  
Objektets rotationsläge  
Menyn Format - Position och storlek... - fliken SnedstÃ¤ll / hÃ¶rnradie  
Menyn Format - Position och storlek... - fliken FÃ¶rklaring  
Snabbmenyn Redigera punkter Snabbmenyn Redigera punkter  
F8 F8  
Ikon på alternativlisten och alternativlisten objektlisten:  
Redigera punkter  
Menyn Format - Teckensnitt (vid ritfunktioner)  
Snabbmenyn Teckensnitt  
Menyn Format - Storlek (vid ritfunktioner)  
Snabbmenyn Storlek  
Menyn Format - Stil (vid ritfunktioner)  
Snabbmenyn Stil  
Menyn Format - Stil - Fet (vid ritfunktioner)  
Snabbmenyn Stil - Fet  
Kommando Ctrl +F  
Ikon på objektlisten:  
Fet  
Menyn Format - Stil - Kursiv (vid ritfunktioner)  
Snabbmenyn Stil - Kursiv  
Kommando Ctrl +K  
Ikon på objektlisten:  
Kursiv  
Menyn Format - Stil - Understrykning (vid ritfunktioner)  
Snabbmenyn Stil - Understrykning  
Kommando Ctrl +U  
Ikon på objektlisten:  
Understruken  
Menyn Format - Stil - Genomstruken (vid ritfunktioner)  
Snabbmenyn Stil - Genomstruken  
Menyn Format - Stil - Skugga (vid ritfunktioner)  
Snabbmenyn Stil - Skugga  
Menyn Format - Stil - Kontur (vid ritfunktioner)  
Snabbmenyn Stil - Kontur  
Menyn Format - Stil - Upphöjt (vid ritfunktioner)  
Snabbmenyn Stil - UpphÃ¶jt  
Kommando Ctrl +H  
Menyn Format - Stil - Nedsänkt (vid ritfunktioner)  
Snabbmenyn Stil - Nedsänkt  
Kommando Ctrl +T  
Menyn Format - Radavstånd (vid ritfunktioner)  
Snabbmenyn Radavstånd  
Menyn Format - Radavstånd - Enradig (vid ritfunktioner)  
Snabbmenyn Radavstånd - Enradig  
Kommando Ctrl +1  
Menyn Format - Radavstånd - 1.5 radig (vid ritfunktioner)  
Snabbmenyn Radavstånd - 1.5 radig  
Kommando Ctrl +5  
Menyn Format - Radavstånd - 2-radig (vid ritfunktioner)  
Snabbmenyn Radavstånd - 2-radig  
Kommando Ctrl +2  
Menyn Format - Justering - Vänster (vid ritfunktioner)  
SnabbmenynJustering - Vänster  
Kommando Ctrl +L  
Ikon på objektlisten:  
Vänsterjusterad  
Menyn Format - Justering - Höger (vid ritfunktioner)  
Snabbmenyn Justering - Höger  
Kommando Ctrl +R  
Ikon på objektlisten:  
Högerjusterad  
Menyn Format - Justering - Centrerad (vid ritfunktioner)  
Snabbmenyn Justering - Centrerad  
Kommando Ctrl +E  
Ikon på objektlisten:  
Justering centrerat horisontellt Centrerad  
Menyn Format - Justering - Marginaljusterad (vid ritfunktioner)  
Snabbmenyn Justering - Marginaljusterad  
Kommando Ctrl +B  
Ikon på objektlisten:  
Marginaljustering  
Menyn Format - FontWork (vid markerat text-ritobjekt)  
Menyn Format - Grupp  
Snabbmenyn Grupp  
Menyn Format - Grupp - Gruppera (textdokument, tabelldokument)  
Menyn Ändra - Gruppera (ritning)  
Snabbmenyn Grupp - Gruppera (formulärobjekt)  
Ikon på objektlisten vid formulärutkast:  
Gruppering  
Menyn Format - Grupp - Upphäva (textdokument, tabelldokument, vid markerad grupp)  
Menyn Ändra - Upphäv gruppering (ritning)  
Snabbmenyn Upphäv gruppering  
Ikon på objektlisten vid formulärutkast:  
Upphäv gruppering  
Menyn Format - Grupp - Lämna (textdokument, tabelldokument, vid markerat objekt inom gruppen)  
Menyn Ändra - Lämna gruppering (teckning)  
Snabbmenyn Lämna gruppering  
Ikon på objektlisten vid formulärutkast:  
Lämna gruppering  
Menyn Format - Grupp - Gå in i (textdokument, tabelldokument, vid markerad grupp)  
Menyn Ändra - Gå in i gruppering (teckning)  
Snabbmenyn Gå in i gruppering  
Ikon på objektlisten vid formulärutkast:  
Gå in i gruppering  
Menyn Format  
Menyn Format - Rad - Höjd...  
Snabbmenyn i ett radhuvud i en öppen databastabell - Radhöjd...  
Menyn Format - Kolumn - Bredd...  
Snabbmenyn i ett kolumnhuvud i en öppen databastabell - Kolumnbredd...  
Menyn Format - Cell... - Flik Tal  
Menyn Format - Mallkatalog... - Ändra / Nytt... - Flik Tal  
Menyn Format - Stylist - snabbmeny Ändra / Nytt... - flik Tal  
Snabbmenyn i ett kolumnhuvud i en öppen databastabell - Kolumnformatering... - Register Format  
Menyn Format - Axel - Y-axel... - Flik Tal (diagramdokument)  
Även som den egna dialogrutan Talformat vid: (Tabell i textdokument) - Format - Talformat... och när man klickat på "Ytterligare format... "i dialogrutan Infoga - FÃ¤ltkommando - Andra...  
Menyn Format - Titel - Flik Justering Menyn Format - Cell... - Flik Justering  
Snabbmenyn i ett kolumnhuvud i en öppen databastabell - Kolumnformatering... - Flik Justering  
Snabbmenyn på ett radhuvud i en öppen databastabell - Tabellformatering...  
Snabbmenyn på ett kolumnhuvud i en öppen databastabell - Kolumnformatering...  
Snabbmenyn på ett radhuvud i en öppen databastabell - Radera rader...  
Menyn Ändra - Spegelvänd (%PRODUCTNAME Draw)  
Menyn Format - Grafik... - fliken Grafik  
Snabbmenyn Spegla (presentationsdokument)  
Menyn Ändra - Spegelvänd - Vertikalt (%PRODUCTNAME Draw)  
Menyn Format - Grafik... - Flik Grafik  
Snabbmenyn Spegla - Vertikalt (presentationsdokument)  
Ikon på bildutrullningslisten på verktygslisten grafikobjektlisten:  
Spegelvänd vertikalt  
Menyn Ändra - Spegelvänd - Horisontellt (%PRODUCTNAME Draw)  
Menyn Format - Grafik... - Flik Grafik  
Snabbmenyn Spegla - Horisontellt (presentationsdokument)  
Ikon på bildutrullningslisten på verktygslisten grafikobjektlisten:  
Spegelvänd horisontellt  
Menyn Ändra - Fördelning... (%PRODUCTNAME Draw)  
Snabbmenyn Fördelning... (%PRODUCTNAME Draw)  
Dölja och fixera förankrade fönster  
Alla förankrade fönster har två ikoner vid kanten mot arbetsområdet och med dem kan du styra fönstervyn.  
Med pilsymbolen döljer respektive visar du fönstret.  
Med den andra symbolen växlar du mellan fixerat och ej fixerat läge.  
I ett ej fixerat läge svävar fönstret över arbetsområdet på ett sådant sätt att fönster som ligger under det delvis täcks.  
Om du inte vill att det ska vara så växlar du över till det fixerade läget, där det förankrade fönstret visas bredvid arbetsområdet.  
Om fönstret förankrats vid arbetsområdets vänstra sida visas följande symboler, beroende på vilket läge som ställts in:  
Visa  
Visa fönstret genom att klicka en gång på pilknappen.  
Dölj  
Dölj fönstret genom att klicka en gång på pilknappen.  
Fixera  
Fixera det genom att klicka en gång på den här kommandoknappen.  
Svävande  
Gör det fritt svävande genom att klicka en gång på den här kommandoknappen.  
AutoShow och AutoHide  
Om Du vid ett dolt fönster klickar på den (förankrade) raden till fönstret öppnas det i AutoShow-läge.  
Fönstret stängs igen automatiskt när Du t ex pekar på arbetsområdet med musen (AutoHide).  
Detta beteende är oberoende av om fönstret är fixerat eller fritt svävande.  
Om ett fönster är i AutoShow-läge visas det så länge musen befinner sig över fönstret och inom dess avgränsningar.  
Även fönsterstorleken kan ändras i AutoShow-läget utan att fönstret stängs.  
Om fönstret förlorar fokus stängs det automatiskt.  
Om Du har förankrat flera fönster bredvid varandra eller över varandra är AutoShow - och AutoHide-beteendet i princip detsamma som vid ett enstaka fönster.  
Du kan även ändra storleken på de enskilda fönstren.  
På så sätt kan Du i AutoShow-läge arbeta med två fönster samtidigt.  
I AutoShow-läget kan Du öppna listrutor i fönstren, anropa snabbmenyer, öppna dialoger och sedan stänga dessa igen utan att fönstret samtidigt stängs.  
AutoHide aktiveras först när Du verkligen inte behöver fönstret längre.  
Dra-och-släpp  
När Du drar ett objekt med musen till ett dolt fönsters (förankrade) rand öppnar sig fönstret även i AutoShow-läge.  
Du kan alltid dra och släppa.  
Snabbmeny Gallery  
Lägg till  
Här kan du definiera i vilken form det markerade grafikobjektet ska integreras i dokumentet.  
Kopia  
Det här kommandot sparar det markerade grafikobjektet som kopia direkt i ditt dokument.  
Det finns då inte längre någon som helst koppling till det ursprungliga grafikobjektet.  
Minnesbehovet för ett dokument är större vid en kopia än vid en länk.  
Länk  
Det här kommandot infogar det markerade grafikobjektet som länk.  
Ett länkat grafikobjekt är bara en slags "hänvisning" till ett originalgrafikobjekt.  
Fördelen är att minnesbehovet är mindre än om du infogar ett grafikobjekt som "kopia".  
Bakgrund  
Här bestämmer du hur bakgrundsgrafikobjektet ska förankras.  
Sida  
Med detta kommando förankras grafikobjektet på sidan.  
Stycke  
Om du väljer det här alternativet förankras grafikobjektet vid stycket.  
Förhandsvisning  
Med detta kommando visas det valda grafikobjektet som enda objekt.  
Om den här funktionen har valts finns en bock framför det här kommandot.  
Genom att återigen välja kommandot Förhandsvisning återställer du den ursprungliga vyn.  
Du kan också välja dessa funktioner (förhandsvisning, ej förhandsvisning) genom att dubbelklicka på respektive grafikobjekt eller med mellanslag.  
Namn  
Här kan du ge ett markerat objekt i ett Gallery-tema ett eget namn.  
Temat får inte vara skrivskyddat.  
När du stänger dialogen Ange namn med OK, övertas namnet som du har matat in där.  
Vid objekt som har en länk till en befintlig fil, visas källans sökväg i parentes efter titeln.  
Radera  
Med detta kommando raderar du det markerade grafikobjektet efter att ha svarat på en kontrollfråga.  
Snabbmeny vid Internet-dokument  
Posternas typ och ordningsföljd i snabbmenyn varierar.  
Det beror dels på vilket objekt som är markerat innan du öppnar snabbmenyn, dels på om dokumentet är skrivskyddat eller i redigeringsläge.  
Öppna  
Om dokumentet är skrivskyddat motsvarar det en "normal" klickning på en länk.  
Öppna i nytt fönster  
Det här kommandot aktiverar länken och öppnar dokumentet i ett nytt fönster.  
Kommandot är bara tillgängligt i redigeringsläge.  
Redigera  
Med det här kommandot väljer du redigeringsläget.  
Du kan också välja redigeringsläget genom att klicka på Redigera på funktionslisten.  
Tillbaka  
Med det här kommandot går du tillbaka till föregående webbdokument.  
Du kan välja den här funktionen genom att klicka på ikonen Bläddra bakåt på funktionslisten.  
Framåt  
Med det här kommandot går du en nivå framåt.  
Det går bara att välja det här kommandot om du redan har gått en nivå bakåt.  
Du kan även klicka på ikonen Bläddra framåt på funktionslisten.  
Spara grafik  
Med det här kommandot öppnar du en dialogruta där du kan spara ett markerat grafikobjekt.  
Kopiera länk  
Med det här kommandot kopierar du länken där muspekaren står till urklippet.  
Kopiera grafik  
Det här kommandot kopierar grafikobjektet där muspekaren står till urklippet.  
Ladda grafik  
Om du har stängt av grafiken kan du göra den synlig igen med det här kommandot.  
Stäng av grafik  
Här kan du välja att grafik i dokumentet ska vara "osynlig".  
Då uppdateras skärmbilden fortare än om grafiken är synlig.  
Stäng av PlugIns  
Med det här kommandot kan du stänga av intregrerade plug-ins.  
Du aktiverar plug-ins genom att välja kommandot igen.  
Spara bakgrund...  
Med det här kommandot kan du spara bakgrunden till en webbsida.  
Du kan sedan t.ex. använda den till din egen hemsida.  
När du har valt Spara bakgrund öppnas en dialogruta där du kan spara grafikobjektet i en valfri katalog.  
Snabbmenyn till aktivitetsfönstren i %PRODUCTNAME  
Sida vid sida  
Detta gäller också om Du har dragit och släppt en aktivitet på en annan aktivitet.  
Horisontal  
Om du har aktiverat flera vyer av ett dokument i en aktivitet med kommandot Nytt fönster, kan du visa alla under varandra med kommandot Horisontal.  
Vertikal  
Om du har aktiverat flera vyer för ett dokument i en aktivitet med kommandot Nytt fönster, kan du visa alla bredvid varandra med kommandot Vertikal.  
Flytande aktivitet  
Med denna omkopplare visas den aktuella aktiviteten i ett nytt, eget fönster.  
När Du klickar igen visas den aktuella aktiviteten som en vanlig aktivitet i hela arbetsområdet.  
Aktivitet alltid synlig  
Med detta kommando blir den aktuella aktiviteten alltid synlig.  
Samtidigt som den blir synlig visas den aktuella aktiviteten som en flytande aktivitet i ett eget fönster.  
När Du klickar igen stängs funktionen av.  
Stäng aktivt fönster  
Om detta är det enda fönstret för en aktivitet, stängs hela aktiviteten.  
Stäng aktivitet  
Den aktiva aktiviteten och alla dess fönster stängs.  
Om Du har ändrat något jämfört med den dokumentversion som finns på datamediet får Du en fråga om Du vill spara ändringarna.  
Nytt  
Här skapar du ett nytt %PRODUCTNAME -dokument.  
I undermenyn bestämmer du med vilken %PRODUCTNAME -komponent du vill arbeta.  
Ett enkelt musklick öppnar ett nytt dokument direkt.  
Ett längre musklick öppnar en undermeny där du kan välja dokumenttyp.  
Om du vill öppna ett dokument som kopia av en dokumentmall, så väljer du kommandot Mallar och dokument.  
En dokumentmall innehåller följande delar:  
Formatmallar för enhetlig utformning av dina dokument  
texter, ramar, kommandoknappar osv.  
Ikon  
Namn  
Funktion  
Textdokument  
Skapar ett nytt textdokument.  
Tabelldokument  
Skapar ett nytt tabelldokument.  
Presentation  
Skapar ett nytt presentationsdokument.  
AutoPilot Presentation öppnas automatiskt om Du inte har valt bort denna funktion.  
Teckning  
Skapar ett nytt teckningsdokument.  
HTML-dokument  
Skapar ett nytt HTML-dokument.  
Samlingsdokument  
Skapar ett nytt samlingsdokument.  
Formel  
Skapar ett nytt formeldokument.  
Etiketter  
Öppnar en dialogruta där Du kan skapa nya etiketter.  
Mallen är ett textdokument.  
Visitkort  
Öppnar en dialogruta där Du kan skapa nya visitkort.  
Mallen är ett textdokument.  
Mallar och dokument  
Öppnar dialogrutan Mallar och dokument.  
Samlingsdokument  
I ett samlingsdokument kan du hantera större projekt, som t.ex. böcker, med hjälp av Navigator för samlingsdokument.  
I samlingsdokumentet lägger du in filer för enskilda kapitel i boken och skapar gemensamma förteckningar för alla deldokument.  
Mallar och dokument  
Dialogrutan Mallar och dokument kan ses som en slags kommandocentral för %PRODUCTNAME -dokument.  
Här finns också alla dokumentmallar, de som medföljde %PRODUCTNAME och de som du själv har skapat.  
Du öppnar dialogrutan via Arkiv - Nytt - Mallar och dokument eller via tangentkombinationen Skift+Ctrl+N.  
I Windows räcker det att dubbelklicka på snabbstartikonen för %PRODUCTNAME %PRODUCTVERSION på aktivitetsfältet.  
Kategori  
Klicka på en kategori här.  
Mallarna eller dokumentet som finns i kategorin visas i listrutan i mitten.  
Listruta  
I listrutan i mitten finns mallarna eller dokumenten Om du klickar på ett objekt visas förhandsvisningen eller dokumentegenskaperna till höger.  
Du öppnar ett dokument resp. öppnar ett nytt dokument som baserar på en mall genom att dubbelklicka.  
Tillbaka  
Ett steg tillbaka i listan med steg som du har utfört i den här dialogrutan.  
Upp en nivå  
Till nästa överordnade mapp (bara under arbetskatalogen).  
Skriv ut  
Utskrift av det valda dokumentet eller den valda mallen.  
Förhandsvisning  
Här ser du en förhandsvisning eller dokumentegenskaper.  
Du byter vy med ikonerna Förhandsvisning och Dokumentegenskaper.  
Förhandsvisning  
Här väljer du förhandsvisning av ett dokument.  
Dokumentegenskaper  
Här väljer du vyn för dokumentegenskaper.  
Du kan ange de här egenskaperna i dialogrutan Egenskaper.  
Administrera  
Öppnar dialogrutan Administrera dokumentmallar.  
Redigera  
Öppnar den valda mallen för redigering.  
Öppna  
Öppnar det valda dokumentet resp. ett nytt dokument som baserar på den valda mallen.  
Om du vill kunna använda en egen mall som inte redan finns i {installpath} / user / template {installpath }\user\template -mappen, måste den här mallen först importeras.  
Klicka på kommandoknappen Kommandon.  
Den valda dokumentmallen överförs till standardkatalogen för dokumentmallar.  
De dokumentmallar som är listade i listrutan Mallar i dialogrutan Nytt administreras i mappen {netinstall} / share / template / swedish ;{userinstall} / user / template C:\{installpath}\share\template\swedish;· C:\{installpath }\user\template.  
Under Verktyg - Alternativ... - %PRODUCTNAME - Sökvägar kan du se sökvägarna för dokumentmallarna och ändra dem.  
Om du registrerar flera sökvägar kan t.ex. alla i ett intranät ha tillgång till de gemensamma mallarna (i ...share...) och ändå använda sina lokala privata mallar (i ...user...).  
Etiketter  
Med den här funktionen administrerar och utformar du etiketter.  
Skriv texten till etiketterna manuellt eller välj innehållet i en databas som etikettext.  
Du kan välja att skriva ut på vanliga pappersark eller på särskilda ark eller rullar med gummerade etiketter.  
Du kan välja bland många olika fördefinierade format, ordnade efter etikettillverkare, och du kan dessutom lätt definiera egna format.  
Du kan också skapa nya dokument för etiketter.  
Det finns en ingående beskrivning om hur etiketter skapas här.  
Nytt dokument  
Med den här kommandoknappen skapar %PRODUCTNAME ett nytt dokument med beteckningen Etiketter1.  
Du kan redigera och komplettera etikettpåskriften i dokumentfönstret.  
Dokumentet kan sparas och skrivas ut.  
Etiketter  
Här bestämmer du dig för etikettpåskrift och väljer etikettformat.  
Påskrift  
Här skriver du texten som ska finnas på alla etiketter.  
Påskrift  
I detta flerradstextfält sammanställer Du påskriften.  
Du kan skriva in texten direkt eller infoga ett databasfält där markören står.  
Adress  
Om Du använder gummerade etiketter för Dina adressutskrifter, markerar Du den här kryssrutan.  
Programmet infogar automatiskt adressuppgifterna i fältet Påskrift.  
Uppgifterna i textfältet baseras på uppgifterna i Användardata under Verktyg - Alternativ - %PRODUCTNAME.  
Databas  
Här väljer Du önskad databas.  
Om Du ska skriva ut etiketter med varierande innehåll, t ex för prisuppgifter, bör Du hämta uppgifterna från en databasfil.  
Tabell  
I det här kombinationsfältet visas en lista över alla tabeller i den valda databasen.  
Posterna beror på urvalet i det vänstra kombinationsfältet Databas.  
Databasfält  
Du kan sätta ihop etikettpåskriften av de olika databasfälten i databasen.  
Välj önskat fält i kombinationsfältet.  
Om Du klickar på pilknapparna till vänster om kombinationsfältet, infogas databasfältet i textfältet Påskrift.  
Under Påskrift visas databasfältsnamnet mellan vinkelparenteser vid markörens position.  
Du måste infoga blanksteg mellan enskilda uppgifter manuellt.  
Om Du vill påbörja en ny rad, trycker Du på Retur när markören står i fältet Påskrift.  
Format  
Här väljer Du ett pappersformat med en viss storlek eller anger egna mått.  
Kontinuerlig  
Välj det här alternativfältet vid utskrift på papper i löpande bana.  
Detta är det format som vanligen används av matrisskrivare.  
Ark  
Välj det här alternativfältet när du ska skriva ut på separata ark.  
Detta är det format som vanligen används av bläckstråle - och laserskrivare.  
Märke  
Välj papperstillverkare i listrutan Märke.  
Varje tillverkare har egna beteckningar på sina format.  
Typ  
Välj en typ i den här listan.  
De uppgifter som visas här gäller alltid den tillverkare som anges i fältet Märke.  
Om den typ som du använder inte finns med på listan, kan du ange egna mått via posten "Användare" under fliken Format.  
Information  
Storleken och placeringen av den valda typen visas i nederkanten av området Format.  
Format  
Här anger du det exakta formatet och placeringen av etiketter eller visitkort på sidan.  
På det här sättet kan du också skriva ut ark och papper i löpande bana som du själv har definierat eller som inte är kända för programmet.  
Horis. avstånd  
Här anger Du det avstånd från vänsterkanten på en etikett eller ett visitkort till vänsterkanten på följande etikett (visitkort) på samma höjd.  
Vert. avstånd  
Här anger Du det avstånd från överkanten på en etikett eller ett visitkort till överkanten på en därunder placerad etikett (visitkort).  
Bredd  
Ange här den faktiska bredden på en etikett eller ett visitkort.  
Höjd  
Ange här den faktiska höjden på en etikett eller ett visitkort.  
Vänster marginal  
Här anger Du avståndet från papperets vänsterkant till vänsterkanten på den första etiketten (första visitkortet).  
Övre marginal  
Här anger Du avståndet från papperets överkant till överkanten på den första etiketten (första visitkortet).  
Kolumner  
Här anger Du antalet etiketter eller visitkort som ska stå intill varandra på samma höjd.  
Rader  
Här anger Du antalet etiketter eller visitkort som ska stå under varandra i samma kolumn.  
Spara...  
Via den här kommandoknappen kommer du till dialogrutan Spara etikettformat.  
Spara etikettformat  
Märke  
Välj märke här.  
Typ  
Ange typ här.  
Tillägg  
Här bestämmer du om du bara vill skriva ut en etikett resp. ett visitkort eller en hel sida.  
Om du inte skriver ut direkt utan skapar ett dokument, anger du under den här fliken om hela sidan i det nya dokumentet ska fyllas, eller om bara en etikett eller ett visitkort ska föras in på den angivna kolumn - och radpositionen.  
Du kan också kontrollera skrivarens konfiguration.  
Hela sidan  
Alla etiketter respektive visitkort skrivs alltid ut på ett ark, eller också skapas en hel sida i det nya dokumentet.  
Enstaka etikett  
Om enbart en enskild etikett (eller ett visitkort) ska skrivas ut eller infogas på den tomma sidan, markerar Du det här alternativet.  
Kolumn  
Här anger Du kolumnnumret för etiketten respektive visitkortet.  
Rad  
Här anger Du radnumret för etiketten respektive visitkortet.  
Synkronisera innehåll  
Markera den här kryssrutan om Du vill redigera en etikett eller ett visitkort och alla ytterligare exemplar ska vara exakta kopior av etiketten eller visitkortet.  
Vid synkronisering övertas också ramattribut, t ex inramning eller bakgrundsgrafik.  
Följande kommandoknappar visas på bildskärmen när Du har markerat kryssrutan Synkronisera innehåll och klickar på kommandoknappen Nytt dokument.  
Synkronisera etiketter  
När Du klickar på den här kommandoknappen, kopieras innehållet i den etikett (det visitkort) som Du redigerar till alla andra etiketter (visitkort) på sidan.  
Funktionen gör det lättare att fylla i data, eftersom Du bara behöver skriva samma data en gång.  
Synkronisera etiketter kan inte användas förrän Du har markerat kryssrutan Synkronisera innehåll och därefter klickat på kommandoknappen Nytt dokument.  
Skrivare  
Här visas namnet på den aktuella skrivaren.  
Ställ in...  
Med den här kommandoknappen öppnar du dialogrutan Ställ in skrivare där du kan ställa in t.ex. sidstorlek, orientering och andra alternativ alltefter skrivartyp.  
Visitkort  
Den här funktionen använder du för att administrera och utforma visitkort.  
Du kan antingen skriva ut på tomt papper eller köpa färdigt material som finns i specialaffärer.  
Det finns ett stort antal format från olika tillverkare.  
Du kan också definiera egna format.  
Medium  
Här anger du formatet för visitkortet.  
Välj bland ett stort antal format från olika tillverkare eller definiera egna format.  
Format  
Här väljer du ett pappersformat med en viss storlek eller anger egna mått.  
Kontinuerlig  
Välj det här alternativfältet vid utskrift på papper i löpande bana.  
Detta är det format som vanligen används av matrisskrivare.  
Ark  
Välj det här alternativfältet när du ska skriva ut på separata ark.  
Detta är det format som vanligen används av bläckstråle - och laserskrivare.  
Märke  
Välj papperstillverkare i listrutan Märke.  
Varje tillverkare har egna beteckningar på sina format.  
Typ  
Välj en typ i den här listan.  
De uppgifter som visas här gäller altlid den tillverkare som anges i fältet Märke.  
Om den typ som du använder inte finns med på listan kan du ange egna mått via posten "Användare" under fliken Format.  
Information  
Storleken och placeringen av den valda typen visas i nederkanten av området Format.  
Visitkort  
Här bestämmer du hur dina visitkort ska se ut.  
Innehåll  
I det här området kan du välja ett AutoText-block för ditt visitkort.  
I listan hittar du AutoText-blocken för det område som är inställt under AutoText - område.  
Välj önskat block genom att klicka med musen.  
AutoText - område  
Här ställer du in området vars innehåll ska visas i innehållslistan.  
Privat  
Under den här fliken finns alla personliga data som ska visas på visitkortet.  
Privata data  
Textfälten i det här området innehåller dina privata data.  
De data du skrev in när du installerade programmet har redan angetts automatiskt.  
Du kan ändra eller komplettera dessa data på menyn Verktyg - Alternativ - %PRODUCTNAME - Användardata eller under den här fliken.  
Förnamn  
Här kan Du ange ytterligare en persons förnamn.  
efternamn  
Här skriver Du in den andra persons efternamn.  
initialer 2  
Här skriver Du in den andra persons initialer.  
Land / Delstat  
I det här textfältet anger Du Ditt land.  
Titel / Yrke  
Här anger Du Din yrkesbeteckning.  
Telefon  
I det här textfältet skriver Du in Ditt privata telefonnummer.  
Mobil  
Om Du har tillgång till mobiltelefon anger Du numret i det här fältet.  
Hemsida  
Här kan du skriva in adressen till din privata hemsida.  
Affärsmässig  
Under den här fliken finns alla affärsdata som ska visas på visitkortet.  
Affärsdata  
Textfälten i det här området innehåller dina affärsdata.  
De data du skrev in när du installerade programmet har redan lagts in automatiskt.  
Du kan ändra eller komplettera dessa data på menyn Verktyg - Alternativ - %PRODUCTNAME - Användardata eller under den här fliken.  
Företag rad 2  
På den här raden kan du skriva in fler företagsuppgifter.  
Slogan  
Skriv in företagets slogan här.  
Land / Delstat  
I det här textfältet kan du skriva in det land där företaget finns.  
Telefon  
I det här fältet skriver du in företagets telefonnummer.  
Mobil  
Om du har tillgång till mobiltelefon anger du numret i det här fältet.  
Hemsida  
Här kan fu skriva in adressen till företagets hemsida.  
Öppna  
Det spelar ingen roll om de är %PRODUCTNAME -dokument eller har externa format.  
Under Verktyg - Alternativ - %PRODUCTNAME - Allmänt kan du välja om du vill använda dialogrutor från %PRODUCTNAME eller från ditt operativsystem när du ska öppna och spara dokument.  
Här beskrivs %PRODUCTNAME -dialogrutan.  
Mer information  
När du öppnar en %PRODUCTNAME -fil som innehåller formatmallar så gäller speciella regler som beskrivs längre ned.  
Upp en nivå  
Om du vill gå upp en nivå i mappstrukturen klickar du på ikonen.  
Den lilla gröna trekanten indikerar att du kan öppna en undermeny genom att klicka där och hålla ner musknappen.  
Den här undermenyn visar de överordnade mapparna.  
Skapa ny katalog  
Med den här ikonen skapar du en ny mapp.  
När du har klickat på ikonen kan du ge mappen ett namn.  
Till standardkatalogen  
Här öppnar du en förinställd mapp eller en mapp som är definierad som standardkatalog för den tilltänkta åtgärden.  
Din "arbetskatalog" eller "standardkatalog "definierar du under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar (Arbetskatalog).  
Visningsområde  
Här visas det urval som passar till de aktuella uppgifterna vid Filnamn och Filtyp.  
Du kan ladda något av de visade dokumenten genom att dubbelklicka på det eller genom att markera det och klicka på kommandoknappen Öppna.  
Kommando Ctrl), kan du klicka på kommandoknappen Öppna och öppna alla filerna samtidigt.  
Du sorterar alla filer genom att klicka på ett kolumnhuvud.  
Om du klickar en gång till sorteras filerna i omvänd ordning.  
Radera - på snabbmeny:  
Raderar markerade filer eller mappar efter säkerhetskontroll.  
Byt namn - på snabbmeny:  
Om du väljer det här kommandot kan du byta namn på en markerad fil eller mapp.  
Filnamn  
Du kan även ange informationen som fullständig URL.  
När du skriver in en URL bör du tänka på att den måste börja med file: / / / eller http: / /.  
Om du skriver in en enhetsbokstav med efterföljande kolon i textfältet, så visas enhetens innehåll i urvalsfönstret.  
Du kan begränsa urvalet av filer i visningsområdet om du skriver in delar av filnamnet tillsammans med platshållare (jokertecken).  
Skriv t ex "a*.*" (alltid utan citattecken) om Du bara vill visa de filer som börjar på "a ".  
Om Du bara minns att ett filnamn har tecknet "3" som tredje tecken och filnamnstillägget "txt", så skriver Du "??3*.txt ".  
Sedan visas bara de filer som motsvarar detta mönster.  
Asterisken "*" står för ett valfritt antal tecken, den får dock inte stå i början eftersom den då skulle tolkas som "alla filer ".  
Frågetecknet "?" står för ett enda valfritt tecken.  
Version  
Om det finns olika dokumentversioner till den markerade filen, så visas de här.  
Du kan skapa och administrera versioner av det dokument som för tillfället är öppet med menykommandot Arkiv - Versioner.  
De olika versionerna av ett dokument öppnas skrivskyddade.  
Filtyp  
I det här fältet väljer du med vilket filter dokumentet ska öppnas.  
I visningsområdet visas nu bara de dokument som motsvarar ditt urval.  
Om du vill se alla filer väljer du "Alla filer (*) (*.*)".  
I början av filtypslistan finns grupper för alla textdokument, tabelldokument o.s.v. som %PRODUCTNAME kan öppna. %PRODUCTNAME bedömer detta med hjälp av filnamnstillägget.  
Mer information om import - och exportfilter.  
När du laddar HTML-filer bör du tänka på att det finns flera filter med namnet Webbsida: filtret i området med de andra %PRODUCTNAME Writer-filtren öppnar dokumentet i %PRODUCTNAME Writer.  
Med filtret i området med de andra %PRODUCTNAME Calc-filtren laddas dokumentet i en %PRODUCTNAME Calc-tabell.  
Detta lämpar sig t.ex. för börsdata som finns i tabellform på Internet.  
Öppna  
När du klickar på den här kommandoknappen avslutas dialogrutan och det valda dokumentet laddas.  
Om inget dokument har markerats, har den här kommandoknappen inte någon funktion.  
Infoga  
När du klickar på den här kommandoknappen infogas den markerade filen vid markörens position i det aktuella dokumentet. (Kommandoknappen Öppna heter Infoga om du har öppnat dialogrutan med menykommandot Infoga - Fil.)  
Bara läsning  
Det går inte att redigera och spara det.  
Men du kan spara dokumentet med ett annat namn, eventuellt i en annan mapp, och sedan redigera det.  
Om den här rutan är markerad är menykommandona som kan ändra dokumentet inte aktiva.  
Spela upp  
Om du klickar på den här kommandoknappen spelas den valda ljudfilen upp.  
Om du klickar igen medan filen spelas upp avslutas uppspelningen.  
Detta är en akustisk "förhandsvisning" av den valda ljudfilen.  
Den här kommandoknappen är bara tillgänglig när en effekt tilldelas ett ljud.  
Tips om hur du öppnar dokument med mallar  
När du öppnar ett %PRODUCTNAME -dokument kontrollerar programmet om dokumentet bygger på en dokumentmall som finns i mappen {installpath} / share / template / swedish {installpath}\share\template\swedish eller i {installpath} / user / template {installpath}\user\template (inklusive de underordnade katalogerna till de här mapparna; eller i de mappar som du har registrerat som mallmappar under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar).  
När du öppnar ett dokument som bygger på en dokumentmall som har ändrats, så visas följande dialogruta:  
Ska dina aktuella mallar användas i det här dokumentet? "  
Om du svarar med Ja laddas dokumentet med den dokumentmall som finns i %PRODUCTNAME.  
De formatmallar som används i dokumentet ersätts med formatmallar med samma namn i %PRODUCTNAME.  
I dokumentet registreras denna ändring först när dokumentet sparas.  
Om du klickar på Nej laddas dokumentet så som det har skapats.  
Formatmallarna i dokumentet ändras inte.  
Om det inte finns någon passande dokumentmall på hårddisken, får du en fråga om mallen ska sökas även vid framtida tillfällen.  
Om Du svarar med Ja letar programmet på nytt efter dokumentmallen när dokumentet laddas nästa gång.  
Detta är ett lämpligt svar om Du t ex vet att formatmallen finns på en nätenhet som för tillfället inte är tillgänglig, men som brukar kunna nås.  
Om Du svarar med Nej och sparar dokumentet, så letar programmet inte längre efter dokumentmallen när dokumentet laddas nästa gång.  
Dokumentet är "frikopplat" från sin formatmall.  
Välj sökväg  
I den här dialogrutan väljer du en mapp som sökväg.  
Dialogrutan motsvarar i stor utsträckning dialogrutan Öppna fil.  
Välja ut  
Klicka här för att välja den visade sökvägen.  
Sökväg:  
I det här kombinationsfältet väljer du den önskade sökvägen eller skriver in en sökväg.  
Filterurval  
I den här dialogrutan väljer du ett importfilter.  
Filter  
I den här listrutan väljer du ett importfilter.  
Den här dialogrutan visas när %PRODUCTNAME inte kan bestämma automatiskt med vilket importfilter filen kan öppnas.  
Välj ett importfilter från listan.  
Installera ett importfilter som saknas (med %PRODUCTNAME Setup -programmet).  
Kontrollera om filen har rätt tillägg för filtypen.  
En fil kan t.ex. ha tillägget .doc även om det är en FrameMaker( tm )-fil.  
Stäng  
Med det här menykommandot stänger du det aktuella dokumentet.  
Om dokumentet är nytt, eller om du ändrat ett befintligt dokument, blir du automatiskt tillfrågad om du vill spara dokumentet innan du stänger det.  
Om Du endast har öppnat ett dokument utan att ändra något stängs det direkt utan att Du får någon fråga.  
Observera dock att %PRODUCTNAME bl a registrerar utskriftsdatum för varje textdokument.  
Om Du skriver ut ett dokument räknas det som en ändring av dokumentet.  
Spara dokument  
Med detta kommando sparar du det aktuella dokumentet  
Om du redigerar ett textblock heter kommandot Spara textblock.  
Spara som  
Här sparar du ditt dokument med ett filnamn och en plats.  
Genom att välja en annan filtyp kan du konvertera dokumentet till ett annat filformat.  
Under Verktyg - Alternativ - %PRODUCTNAME - Allmänt kan du välja om du vill använda dialogrutor från %PRODUCTNAME eller från ditt operativsystem när du ska öppna och spara dokument.  
Här beskrivs %PRODUCTNAME -dialogrutan.  
Information som du anger under Arkiv - Egenskaper ändras inte när dokumentet sparas, även om du använder ett nytt namn.  
Eftersom en titel som du anger under Arkiv - Egenskaper - Beskrivning även visas i titellisten i %PRODUCTNAME, bör du ändra sådana poster för att undvika förväxlingar.  
Du ombeds alltid att ange plats och namn.  
Den här filtypen används t.ex. till datorns konfigurations - och startfiler.  
Om du har öppnat en HTML-källtext heter kommandot Exportera källtext Om det rör sig om tecknings - och presentationsdokument och du väljer kommandot Exportera heter den här dialogrutan Exportera.  
Upp en nivå  
Om du vill gå upp en nivå i katalogstrukturen klickar du på ikonen Upp en nivå.  
Den lilla gröna triangeln signalerar att du med en lång klickning kan öppna en undermeny.  
Den här menyn visar respektive överordnad katalog.  
Här kan du välja en katalog.  
Skapa ny katalog  
Med den här ikonen skapar du en ny mapp.  
När du har klickat på ikonen kan du skriva ett namn för mappen.  
Till standardkatalogen  
Här öppnar du en katalog som redan har ställts in resp. en katalog som har definierats som standardkatalog för den här åtgärden.  
Visningsområde  
Här visas ett filurval enligt inställningen av Filtyp som du har gjort.  
Filnamn  
I det här kombinationsfältet kan du skriva namnet på dokumentet som ska sparas direkt.  
Du kan också ange namnet som en fullständig URL-adress.  
Filtyp  
I det här kombinationsfältet bestämmer du formatet på det dokument som ska sparas.  
I visningsområdet syns bara de dokument som motsvarar de val som du har gjort här.  
Mer information om filtyper finns i avsnittet Information om import - och exportfilter.  
Se därför alltid till att först spara dokumentet i %PRODUCTNAME -programmets format innan du exporterar det till externa format.  
Om du vill kunna öppna och redigera filen i en äldre version av %PRODUCTNAME, måste du spara den i motsvarande format (t.ex. %PRODUCTNAME Writer 2.0).  
Spara  
Med den här kommandoknappen stänger du dialogrutan och sparar dokumentet med det angivna namnet.  
Om du har angett ett namn på ett dokument som redan finns, ber %PRODUCTNAME dig att först bekräfta att dokumentet ska skrivas över.  
Antingen bekräftar du det - då ersätter det nya dokumentet det gamla - eller också avbryter du genom att klicka på kommandoknappen Avbryt.  
Spara med lösenord  
Genom att markera den här rutan förhindrar du att obehöriga läser eller ändrar ditt dokument.  
Innan skyddet träder i kraft visas dialogrutan Mata in lösenord där du anger och bekräftar ditt lösenord.  
Spara med lösenord är bara möjligt för de XML-baserade dokumentformaten från %PRODUCTNAME %PRODUCTVERSION.  
Automatiskt filnamnstillägg  
Om du har markerat den här rutan, sparas filen med det filnamnstillägg som motsvarar den filtyp som du har valt.  
Redigera filterinställningar  
Öppnar dialogrutan Textexport för filtypen "Text CSV".  
Markering Markering  
Du markerar den här rutan om du bara vill exportera markerade objekt från %PRODUCTNAME Draw till ett externt grafikformat.  
Om den här rutan inte är markerad, exporteras hela sidan.  
För filtypen Webbsida exporteras alltid hela sidan.  
Du markerar den här rutan om du bara vill exportera de markerade elementen från %PRODUCTNAME Impress till ett externt grafikformat.  
Om den här rutan inte är markerad, exporteras hela sidan.  
För filtypen Webbsida exporteras alltid hela sidan.  
Egenskaper för  
Här hittar du allmän information om det aktuella dokumentet.  
Du kan alltså alltefter tillämpning se t.ex. antalet ord och tecken i texten eller det datum då dokumentet skapades.  
Du kan också själv ange egenskaper och ändra dem, t.ex nyckelord eller ett namn som inte hör ihop med filnamnet.  
Du kan också definiera nya fält med ytterligare textinformation.  
Om dokumentet är skrivskyddat, är även alla egenskapsfält skrivskyddade. (Du kan placera markören i fälten men inte ändra innehållet.)  
Annars övertas de i den nya filen, vilket kan leda till förväxlingar.  
Med kommandot Egenskaper... kan du även tillfoga kompletterande information till dokumentet.  
Vidare finns det en statistikfunktion som ger information om dokumentinnehåll och lagringsdata.  
Dessutom finns det en statistikfunktion som ger information om dokumentinnehållet.  
Vid delningskonflikter eller om du saknar behörighet till ett dokument har du inte tillgång till funktionerna under de enskilda flikarna.  
Då kan du bara läsa dokumentinformationen under några av flikarna.  
Du ser följande flikar:  
Beskrivning  
Den här fliken använder du när du ska ange information om dokumentet.  
HTML-import och export  
När dokumentet sparas som HTML-fil, exporteras fältens innehåll automatiskt som följande META NAME -taggar.  
Du använder den här funktionen till att föra in t.ex. upphovsrättsinformation eller nyckelord för de automatiska sökmotorerna på din sida, även om orden inte förekommer i läsbar text på sidan.  
Rubrik  
<TITLE>  
Tema  
<META NAME=" CLASSIFICATION "CONTENT="fältinnehåll ">  
Nyckelord  
<META NAME=" KEYWORDS "CONTENT="fältinnehåll ">  
Beskrivning  
<META NAME=" DESCRIPTION "CONTENT="fältinnehåll ">  
Informationsfält 0...3  
<META NAME=" informationsfältnamn "CONTENT="fältinnehåll ">  
Importanvisningar  
Ytterligare META-taggar som vid import automatiskt utvärderas i %PRODUCTNAME är <META HTTP-EQUIV=" REFRESH"...> och <META NAME="... "...> där NAME är AUTHOR, CREATED, CHANGED, CHANGEDBY, DESCRIPTION, KEYWORDS eller CLASSIFICATION.  
Dessutom förs de första fyra META-taggarna med NAME-alternativ in som användaregenskaper i dokumentet.  
När du importerar HTML-taggar kan du ange i dialogrutan Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet om okända taggar ska importeras som fält eller hoppas över.  
Till de kända taggarna hör META-taggarna när de hänvisar till ett HTTP-EQUIV - eller NAME-alternativ.  
I så fall används uppgiften i det alternativet medan övriga alternativ hoppas över.  
Undantag: en <META NAME=" GENERATOR "...> hoppas genomgående över.  
Om dessa kända taggar inte hoppas över, importeras de som anteckningar.  
De blir i stället (liksom kommentarer och META-taggar) infogade i den första tabellcellen.  
Kommentarer, META-taggar och skript som står omedelbart före ett sidhuvud, infogas inte i detta utan förblir förankrade i huvuddokumentet.  
Alla kommentarer, META-taggar och skript som finns i HEAD-avsnittet förankras på detta sätt till dokumentets första stycke och exporteras senare tillbaka till HEAD.  
Exportinformation  
Vid export i HTML exporteras en anteckning som börjar med "<META" och slutar med "> "inte som en kommentar utan i sin helhet som META-tagg.  
Anteckningar och skript-fält som står i början av det första stycket i ett dokument (men inte i sidhuvudet) exporteras i HTML-dokumentets HEAD-avsnitt.  
Om dokumentet börjar med en tabell, betraktas det första stycket i den första tabellcellen.  
Rubrik  
I det här textfältet anger Du dokumentets rubrik.  
Den visas på rubrikraden.  
Tema  
I det här textfältet anger Du dokumentets ämne.  
Nyckelord  
I det här textfältet anger Du olika nyckelord för dokumentet.  
Beskrivning  
Här ger Du en beskrivning av dokumentet.  
Allmänt  
Under fliken Allmänt finns allmän information om det aktuella dokumentet, t.ex. sökväg till mappen, vilken mall som används, datum då dokumentet skapats och ändrats, författare etc.  
Fil  
Här visas filnamnet och filikonen.  
Om filnamnet är längre än textfältet visas början på filnamnet.  
Typ:  
Här visas information om det aktuella dokumentets filtyp.  
Plats:  
Här anges var det laddade dokumentet är placerat.  
Storlek:  
Här visas storleken för det aktuella dokumentet i byte.  
Skapat:  
Här visas datum och klockslag när första versionen av dokumentet sparades.  
Om Du öppnar ett dokument i rent textformat skapar %PRODUCTNAME ett %PRODUCTNAME Writer-textdokument av det och visar det på bildskärmen.  
Du kan utföra alla typer av formatering som är tillgängliga för %PRODUCTNAME Writer-textdokument, även formatering som inte kan visas i rena textfiler.  
Detta visar att dokumentet på bildskärmen är något mer (eller något annat) än ursprungsdokumentet som kanske bara finns i rent ASCII-format.  
Det dokument Du ser är ju faktiskt ett nytt dokument!  
När Du sedan sparar kan Du bestämma om Du vill spara som ett rent textdokument utan formatering eller som ett %PRODUCTNAME Writer-textdokument.  
Ändrat:  
Här visas datum och klockslag när dokumentet senast ändrades.  
Version:  
Här anges dokumentets versionsnummer.  
Detta tilldelas automatiskt varje gång som du sparar dokumentet.  
Utskrivet:  
Datum och klockslag för senast utskrift visas här.  
Mall:  
Om du har använt en dokumentmall visas dokumentmallens namn här.  
Redigeringstid:  
I det här fältet visas total redigeringstid för dokumentet.  
Den totala tidsåtgången fram till det tillfälle då dokumentet senast sparats visas.  
Den totala redigeringstiden registreras i dokumentets egenskaper varje gång som Du sparar filen.  
Skrivskyddad  
Den här kryssrutan visas bara när du öppnar den här fliken med kommandot Egenskaper på snabbmenyn för ett oöppnat dokument.  
Om du markerar den här rutan förser du det oöppnade dokumentet med attributet "skrivskyddat".  
Då kan det bara öppnas för läsning.  
Ett oöppnat dokument kan vara skrivskyddat utan att ha attributet "skrivskyddad".  
Det kan t.ex. vara fallet om en annan användare redan har öppnat dokumentet.  
Använd användardata  
Om den här rutan är markerad sparas användarens namn tillsammans med dokumentet.  
Namnet visas under Arkiv - Egenskaper - Allmänt.  
Radera  
Med den här kommandoknappen ändrar Du skapandedatum till aktuellt datum och författarens namn till den aktuella användarens namn.  
Värdena för Ändrat och Utskrivet raderas.  
Redigeringstid ställs på 0 och versionsnumret ställs på 1.  
Användare  
Här kan du ange fyra valfria uppgifter om dokumentet.  
Info 0 till Info 3  
I de här textfälten kan du föra in valfri information.  
Infofält...  
Genom att klicka på den här kommandoknappen öppnar Du en dialogruta där Du kan ange namn på de olika infofälten.  
Redigera informationsnamn  
I den här dialogrutan kan Du ändra informationsnamnen.  
Namn  
I det här området i dialogrutan finns de inmatningsfält där du kan ange namn för de olika infofälten i dokumentet.  
I de fyra textfälten skriver Du rubrikerna på infofälten 0 till 3.  
Om Du bekräftar med OK, visas uppgifterna i användarregistret.  
Statistik  
Under fliken Statistik hittar du statistiska uppgifter om det aktuella dokumentet: antal sidor vid utskrift, antal tabeller, grafiska objekt och OLE-objekt i dokumentet, antal stycken, ord och tecken. och celler.  
Antal sidor:  
Här hittar du det totala antalet sidor när dokumentet skrivs ut.  
Tabellantal; dokumentAntal tabeller:  
Här anges det totala antalet tabeller som finns i dokumentet.  
Tabeller som infogats som OLE räknas inte med.  
Antal celler:  
Här visas antalet icke-tomma celler i tabellerna.  
Antal grafikobjekt:  
Här visas det totala antalet grafiska objekt som finns i dokumentet.  
I beräkningen ingår både de grafiska objekt som sparats i dokumentet och sådana som det finns en referens till.  
Grafiska objekt som infogats som OLE räknas inte med (se menyn Infoga - Grafik).  
Antal OLE-objekt:  
Här visas det totala antalet OLE-objekt som finns i dokumentet, inklusive tabeller och grafiska objekt som infogats som OLE.  
Antal stycken:  
Här visas det totala antalet stycken i dokumentet.  
Även tomma stycken räknas med.  
Antal ord:  
Här visas det totala antalet ord i dokumentet.  
Det minsta ord som räknas är exakt ett tecken långt.  
Avgränsare  
I detta fält kan Du ange de tecken som ska fungera som avgränsare vid beräkningen.  
Vanligtvis betraktas ord som ett enda ord om de t ex binds samman med tecknet /.  
Om Du vill att ord som är sammanfogade på detta sätt ska räknas vart för sig, så anger Du det önskade tecknet i inmatningsfältet för avgränsare.  
Detta gör att t ex Persson / Schyman eller Persson&Schyman räknas som två ord vid beräkningen.  
Du kan ange vilka tecken som helst.  
Specialtecken och icke utskrivbara tecken kan även anges hexadecimalt.  
För ett tecken enligt ASCII -Code 255 skriver Du \xff (x[hexadecimalt tal]).  
Specialtecken som \n (LineFeed) och \t (Tab) stöds också.  
Antal tecken:  
Här hittar du det totala antalet tecken i dokumentet inklusive alla mellanslag.  
Kontrolltecken, t.ex. stycketecken, räknas inte.  
Antal rader:  
Här visas det totala antalet rader i dokumentet.  
Uppdatera  
Om du klickar på den här kommandoknappen beräknas och visas antalet rader i dokumentet.  
Internet  
Under fliken Internet bestämmer du om ett laddat HTML-dokument ska ladda ett annat HTML-dokument efter en viss tid som går att ställa in.  
Här bestämmer Du om och efter hur lång tid ett följande dokument till det aktuella dokumentet ska laddas.  
Genom att på detta sätt "länka" flera dokument till varandra kan Du t.ex. skapa självgående presentationer.  
Men Du kan också låta ladda om samma dokument gång på gång, om det t.ex. innehåller länkar till databaser vars innehåll hela tiden kan ändras.  
Ladda automatiskt efter  
Markera det här fältet om det följande dokumentet ska laddas automatiskt efter det antal sekunder som anges i rotationsfältet Sekunder.  
Sekunder  
I det här rotationsfältet anger Du efter hur lång tid laddningen av det följande dokumentet ska ske.  
URL  
Ange här fullständig URL till det följande dokumentet.  
Ram  
Här anger Du de målramar som används som standard för alla hyperlänkar i det aktuella dokumentet, om inte en annan målram är definierad i själva hyperlänken.  
Du kan även välja bland standardvärdena i listan till höger som öppnas om Du klickar på knappen med nedåtpilen.  
Standardvärdena har följande innebörder:  
Standard  
Betydelse  
Förinställda målramstyper  
Val bland de ramar i dokumentet som redan har fått namn  
_self  
Det följande dokumentet visas i samma ram  
_blank  
Det följande dokumentet visas i en tom, ny ram  
_parent  
Om det inte finns någon, visas dokumentet i samma ram.  
_top  
Om det inte finns någon, visas dokumentet i samma ram.  
Dokumentmall  
Du kan även spara det aktuella dokumentet som dokumentmall.  
Adressbokskälla  
Administrera  
Öppna dialogrutan Administrera dokumentmallar där du kan kopiera, radera, redigera, importera och exportera dokumentmallar och skapa nya dokumentmallar.  
Här definierar du även standardmallar.  
Vänster och höger listruta (dokumentmallar / dokument)  
I den undre listrutan väljer du om dokumentmallar eller dokument ska visas.  
Här visas motsvarande filer.  
Välj om dokumentmallar ska listas i urvalslistrutan i listrutan Dokumentmallar.  
Välj Dokument om dokumentfiler ska visas i listrutan ovanför.  
Vid visningen av dokumentmallar visas de mappar och dokumentmallar som finns i sökvägen för dokumentmallar, samt deras innehåll, i listrutan.  
Mappsymbolerna representerar då de olika mallkategorierna.  
Dokumentmallarna sparas som standard i template-mappen i Office-katalogen: färdiga dokumentmallar i {installpath} / share / template / swedish {installpath}\share\template\swedish och egna dokumentmallar i {installpath} / user / template {installpath }\user\template.  
Den här inställningen gör du under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar.  
Om du sedan dubbelklickar på en dokumentmalls ikon visas ikonerna Mallar och Konfiguration.  
Om du dubbelklickar på mallsymbolen listas alla formatmallar som används i dokumentet enskilt, t.ex. stycke - och teckenformatmallar.  
Om du dubbelklickar på konfigurationssymbolen visas de olika konfigurationerna, i den mån du har definierat egna konfigurationer för dokumentet i dialogrutan Anpassa.  
Om du visar dokumentmallarna i en listruta och dokumenten i den andra listrutan kan du dra-och-släppa de enskilda formatmallarna eller konfigurationerna från ett dokument till en dokumentmall (och vice versa).  
Välj formatmall eller konfiguration och dra den med musen till dokumentposten.  
Om det redan finns en formatmall av samma typ och med samma namn i ett dokument får du en kontrollfråga om den befintliga formatmallen ska ersättas.  
Kommandon  
Om du klickar på den här kommandoknappen får du tillgång till olika kommandon för hantering av dokumentmallarna.  
Vilka av de kommandona i undermenyn som är tillgängliga beror på den aktuella markeringen (dokument, dokumentmall eller dokumentmallsmapp).  
I undermenyn finns följande kommandon:  
Nytt  
På det här sättet skapar du ett nytt mallområde (mapp).  
Standardbeteckningen "namnlös" är markerad.  
Klicka sedan utanför namnet i listrutan.  
Radera  
Med det här kommandot tas det mallområde som är markerat i listrutan eller den markerade dokumentmallen bort.  
Innan raderingen genomförs får du en kontrollfråga.  
Redigera  
Med det här kommandot laddar du dokumentmallen som är markerad i listrutan.  
Importera mall  
Sedan väljer du Importera mall.  
Då visas en standarddialog där du kan välja en dokumentmall (se dialogrutan Öppna).  
Förinställningen är att katalogen som är angiven som "Arbetskatalog" (se Verktyg - Alternativ - %PRODUCTNAME - Sökvägar) öppnas.  
Exportera mall  
Med det här kommandot kan du exportera mallen som är markerad i listrutan.  
Mallen sparas med ett nytt namn.  
En standarddialogruta visas där dokumentmallar kan sparas (se dialogrutan Spara som).  
Förinställningen är att katalogen som är angiven som "Arbetskatalog" öppnas (se Verktyg - Alternativ - %PRODUCTNAME - Sökvägar).  
Skriv ut  
Om du vill skriva ut inställningarna i formatmallarna dubbelklickar du på dokumentmallen i listrutan, väljer Mallar och öppnar snabbmenyn.  
Välj sedan Skriv ut.  
Skrivarinställningar...  
Innan du skriver ut kan du göra skrivarinställningar här.  
Standarddialogrutan där du kan välja skrivare visas.  
Du kan välja en annan skrivare eller ändra inställningarna för den aktuella skrivaren.  
Uppdatera  
Visningen i listrutorna uppdateras.  
Definiera som standardmall  
Med det här kommandot definierar du det malldokument, som är markerat i dialogrutan, som standardmall för alla nya dokument av den här typen.  
Återställ standardmall  
Här öppnas en undermeny där alla dokumenttyper visas som har definierats som standardmallar.  
Välj den typ för vilken den ursprungliga förinställningen ska gälla.  
Adressbok  
Här öppnar du dialogen Mallar: adressbokstilldelning.  
Fil...  
Om du vill kopiera mallar eller konfigurationer från ett %PRODUCTNAME -dokument markerar du dokumentet i listrutan och väljer Fil.  
Då visas en standarddialogruta där du kan välja fil (se dialogrutan Öppna).  
Det dokument som är markerat där visas i listrutan.  
Mallar: adressbokstilldelning  
Här väljer du vilken tabell från vilken datakälla som ska användas som adressbok i %PRODUCTNAME.  
Adressbokskälla  
Välj datakälla och tabell för adressboken.  
Datakälla  
Välj datakällan för adressboken här.  
Tabell  
Välj tabellen för adressboken här.  
Administrera  
Här öppnar du dialogen Administrera datakällor.  
Fälttilldelning  
Bestäm fälttilldelningen för adressboken här.  
(Fältnamn)  
Välj ut den post i kombinationsfältet som motsvarar %PRODUCTNAME -adressboksfältet.  
Efter "Företag" väljer du t.ex. datafältet som motsvarar %PRODUCTNAME -adressboksfältet "Företag "i din adressbok.  
Spara (dokumentmallar)  
Här sparar du det aktuella dokumentet som ny dokumentmall.  
Den här funktionen gör att du senare kan öppna ett nytt dokument som ser ut exakt som det du sparat som dokumentmall.  
Ny dokumentmall  
Här anger du namnet på den dokumentmall som ska sparas.  
Mallar  
Här bestämmmer du i vilken kategori din nya dokumentmall arkiveras.  
Kategorier  
Här väljer du en kategori som den nya dokumentmallen ska sparas i.  
Om du vill skapa en ny kategori, klickar du på kommandoknappen Administrera....  
Mallar  
I den här listrutan visas de dokumentmallar som finns i den markerade kategorin.  
Redigera  
Om du klickar på den här kommandoknappen laddas dokumentmallen som är markerad i mallområdet för redigering.  
Administrera...  
Med kommandoknappen Administrera... öppnar du dialogrutan Administrera dokumentmallar.  
Redigera  
Här öppnar du en dialogruta där du kan öppna en dokumentmall.  
Den motsvarar dialogrutan Öppna.  
Förhandsgranskning / sidutskrift FÃ¶rhandsgranskning  
Här aktiverar och deaktiverar du förhandsgranskningen av dokumentet.  
På det sättet kontrollerar du redan före utskriften hur t.ex. sidindelningen ser ut.  
Förhandsgranskningslisten innehåller bl.a. ikoner för bläddring i flersidiga dokument eller för samtidig visning av flera sidor (se beskrivningen av förhandsgranskningslisten listen "Förhandsgranskning ").  
Bläddra genom vyn med Ctrl + Page Up och Ctrl + Page Down.  
I förhandsgranskningen kan du inte göra några ändringar i dokumentet.  
Om du dubbelklickar på ett ställe i förhandsgranskningen aktiveras dokumentets normalvy igen.  
Använd även förhandsgranskningen till att skriva ut flera dokumentsidor på en papperssida.  
I %PRODUCTNAME Writer hittar du ikonen Utskriftsalternativ på listen "Förhandsgranskning".  
Om du klickar på ikonen öppnas en dialogruta där du kan välja inställningar för utskrift av flera sidor.  
Skriv ut  
Med menykommandot Skriv ut kan du definiera olika utskriftsalternativ och skriva ut det aktuella dokumentet.  
Skrivare  
Du kan också välja att skriva ut till en fil.  
Namn  
I den här listrutan väljer du vilken av de installerade skrivarna du vill använda.  
Status  
Här visas om skrivaren är redo och om det rör sig om standardskrivaren.  
Typ  
I det här textfältet visas namnet på den använda skrivardrivrutinen.  
Plats  
Här anges skrivarporten.  
Kommentar  
Om du eller skrivarens tillverkare har försett skrivardrivrutinen med en kommentar, så visas den här.  
Egenskaper  
Den här kommandoknappen öppnar en dialogruta där du kan ställa in skrivarens egenskaper.  
Den här dialogrutan tillhandahålls av skrivardrivrutinen, därför ser dialogrutan olika ut beroende på vilken skrivare som används.  
Detaljerad information hittar du i dokumentationen för skrivaren.  
Skriv ut till fil  
Markera här om du vill skriva ut direkt till en fil.  
...  
Den här kommandoknappen öppnar dialogrutan Spara som där du kan välja mapp och eventuellt det filnamn till vilket du vill skriva ut.  
Utskriftsområde  
Här väljer du vilka av dokumentets sidor som ska skrivas ut.  
Om du har definierat ett utskriftsområde i %PRODUCTNAME Calc, skrivs bara utskriftsområdet ut.  
Allt  
Välj det här alternativet om du vill att alla sidor i det aktuella dokumentet ska skrivas ut.  
Sidor  
Bara de sidor som anges i textfältet skrivs ut.  
Om du vill skriva ut enstaka sidor, skiljer du sidnumren åt med semikolon:  
3; 8; 10.  
3-12.  
Om sidorna 3, 6 och 9 till 14 ska skrivas ut, anger du:  
3; 6; 9-14.  
Markering  
Bara de markerade texterna eller objekten i dokumentet skrivs ut.  
Kopior  
Här anger du hur många exemplar som ska skrivas ut.  
Exemplar  
I det här rotationsfältet anger du hur många exemplar som ska skrivas ut totalt.  
Sortera  
Markera den här rutan om exemplaren ska skrivas ut sammanhängande, d.v.s. först det första exemplaret komplett, sedan det andra osv.  
Om inte alla de celler finns med på utskriften som Du anser borde skrivas ut, så kan Du kontrollera om Du har definierat ett utskriftsområde.  
Ifall ett sådant finns definierat, så skrivs bara utskriftsområdets innehåll ut!  
Fler  
Om du klickar på den här kommandoknappen visas dialogrutan Skrivaralternativ.  
Om du klickar på den här kommandoknappen visas dialogrutan Skrivaralternativ.  
Dialogrutan motsvaras av en sida i alternativdialogen som du öppnar genom att välja Verktyg - Alternativ - Textdokument - Skriv ut.  
Här ställer du in vilken information som inte ska finnas med på utskriften, hur anteckningarna ska behandlas vid utskriften, vilket pappersmagasin som ska användas med mera.  
Inställningarna i dialogrutan Skrivaralternativ gäller bara för det aktuella dokumentet.  
Om du vill använda enskilda inställningar i denna dialogruta generellt för alla andra dokument, kan du under Verktyg - Alternativ - Textdokument - Skriv ut definiera dem som globala inställningar för alla dokument av detta slag i %PRODUCTNAME.  
Via kommandoknappen Fler kommer du till dialogrutan Skrivaralternativ.  
Den här dialogrutan motsvaras av en sida i alternativdialogen som du öppnar genom att välja Verktyg - Alternativ - Tabelldokument - Skriv ut.  
Via kommandoknappen Fler kommer du till dialogrutan Skrivaralternativ.  
Den här dialogrutan motsvaras av en sida i alternativdialogen som du öppnar genom att välja Verktyg - Alternativ - Teckning - Skriv ut.  
Via kommandoknappen Fler kommer du till dialogrutan Skrivaralternativ.  
Den här dialogrutan motsvaras av en sida i alternativdialogen som du öppnar genom att välja Verktyg - Alternativ - Teckning - Skriv ut.  
Om du klickar på den här kommandoknappen visas dialogrutan Skrivaralternativ som motsvarar dialogrutan Inställningar under Verktyg - Alternativ - Formel.  
I den senare dialogrutan gör du inställningar som gäller för alla dokument, medan inställningarna i dialogrutan Skrivaralternativ bara gäller för den aktuella utskriften.  
Under Unix visas Windows-specialtecknen 128 - 160 vid utskrift.  
Detta gör att det är möjligt att skriva ut ett dokument, som har skapats med %PRODUCTNAME för Windows och som t.ex. innehåller typografiska tecken, på en PostScript-skrivare under Unix.  
Specialtecknen syns bara på utskriften - eftersom Xservern inte känner till dem, visas de inte på bildskärmen.  
FontMetric (teckenbredd) stämmer bara exakt för Monospaced Fonts, för andra teckensnitt är den ungefärlig.  
Genom Environment-variabeln STAR_SPOOL_DIR kan du ange en katalog där spoolfiler för skrivaren X ska placeras under Unix.  
Exempel:  
setenv STAR_SPOOL_DIR / usr / local / tmp (i csh / tcsh) eller  
export STAR_SPOOL_DIR= / usr / local / tmp (i sh / bash)  
I konfigurationsprogrammet spadmin kan du göra den här och andra inställningar i en dialogruta.  
Öppna dialogrutan Koppla.  
Inställningarna för kön kan du även definiera som allmänna förinställningar genom att klicka på en kommandoknapp.  
Ställ in skrivare  
Med det här kommandot öppnar du en dialogruta med information om skrivaren.  
Du kan också ändra egenskaperna om du går till dialogrutan för den enskilda skrivaren.  
Som regel kan du t.ex. välja pappersstorlek och pappersmagasin i skrivarens dialogruta.  
Detta förutsätter att Du har angett att ett sådant meddelande ska skickas (t ex i %PRODUCTNAME Math).  
Eftersom det kan dröja lite innan ett sådant meddelande laddas, visas ibland en förloppsindikator med meddelandet "Anpassa objekt...".  
Skrivare  
I detta område finns uppgifter från skrivardrivrutinen.  
Beroende på skrivare kan Du göra olika inställningar.  
Namn  
Du kan också välja en annan installerad skrivare.  
Om Du redan har skrivit ut Ditt dokument står namnet på den senast använda skrivaren i denna listruta.  
Om Du har flera skrivardrivrutiner installerade på datorn kan Du välja en av dem i listrutan.  
Status  
Här visas om skrivaren är driftklar och om det är standardskrivaren.  
Typ  
I detta textfält finns namnet på den skrivardrivrutin som används.  
Plats  
Här visas skrivaranslutningen.  
Kommentar  
Om Du eller skrivartillverkaren har försett skrivardrivrutinen med en kommentar så visas den här.  
Egenskaper...  
Om du klickar på den här kommandoknappen öppnas dialogrutan Egenskaper för skrivardrivrutinen.  
Eftersom den här dialogrutan kommer från skrivartillverkaren är den utformad på olika sätt beroende på vilken skrivare som används.  
Tänk på att sidorienteringen stående eller liggande format som du kan ställa in i skrivaregenskaperna, måste stämma överens med det sidformat som du har ställt in med hjälp av Format - Sida.  
Du måste alltid installera en standardskrivare i systemet för att dokumenten i %PRODUCTNAME ska kunna visas på bildskärmen så som de ser ut vid utskrift.  
I Windows installerar du en standardskrivare via Start-menyn - Inställning - Kontrollpanelen - Skrivare.  
I Unix använder du programmet spadmin när du ska registrera en standardskrivare för %PRODUCTNAME.  
Skicka  
Med det här kommandot öppnar du en undermeny med kommandon för att skicka det aktuella dokumentet som e-post.  
Om det aktuella dokumentet är ett textdokument, innehåller undermenyn ytterligare några kommandon.  
Du kan överföra dispositionen till ett %PRODUCTNAME Impress-dokument eller till urklippet, skapa ett AutoUtdrag, ett samlingsdokument eller ett HTML-dokument.  
Dokument som e-post  
Skapa samlingsdokument  
Skapa HTML-dokument  
Skapa AutoUtdrag...  
Skicka dokument som e-post  
Med det här kommandot skickar du det aktuella dokumentet som e-post.  
Kommandot öppnar det program som är registrerat som standard-e-postprogram i systemet.  
Det aktuella dokumentet är redan infogat som e-postbilaga där.  
Samlingsdokumentets namn och sökväg  
Här skapar du ett samlingsdokument utifrån ett textdokument.  
För varje kapitel, som börjar med en styckeformatmall som du har valt, sparas automatiskt ett nytt deldokument.  
När du har valt kommandot öppnas dialogrutan Samlingsdokumentets namn och sökväg där du anger namn och sökväg för det samlingsdokument som ska skapas.  
Dialogrutans funktion motsvarar dialogrutan Spara fil.  
Samlingsdokumentet får automatiskt filnamnstillägget .sxg (t.ex. "Samling.sxg").  
Deldokumentens namn baseras på detta.  
Det första deldokumentet får samma namn som samlingsdokumentet med tillägget 1, men med filnamnstillägget .sxw ("Samling1.sxw").  
Det andra deldokumentet får namnet "Samling2.sxw" och så vidare.  
Där visas namnen på de deldokument som du har skapat.  
Dubbelklicka på ett namn eller markera det och klicka på Redigera i Navigator om du vill redigera ett deldokument.  
Visningsområde  
Filnamn  
Aktuell mall  
Välj styckeformatet som ska fungera som avgränsning.  
I normala fall delar du utgångsdokumentet vid de stycken som har formaterats med formatet "Överskrift 1".  
På så vis blir varje kapitel till ett eget deldokument.  
Här kan du också välja en annan mall bland styckeformatmallarna som används i dokumentet.  
Filtyp  
Spara  
Automatiskt filnamnstillägg  
Avsluta  
Med det här kommandot avslutar du %PRODUCTNAME och alla öppna dokument.  
Du blir tillfrågad om du vill spara ändringarna.  
Om du har startat en s.k. referensdialog, t.ex. funktionsautopiloten i %PRODUCTNAME Calc, måste du stänga den innan du kan avsluta %PRODUCTNAME.  
Spara allt  
Med det här kommandot sparar du alla öppna dokument.  
Denna funktion kan du bara använda om du redigerar minst två dokument.  
Dokumenten sparas med aktuella sökvägar och namn och de gamla versionerna skrivs över.  
Där anger Du namn på filen och var den ska sparas.  
Versioner  
Här kan du spara flera versioner av ett dokument.  
Du kan spara en ytterligare version av ett dokument med kommandot Versioner.  
I dialogrutan Versioner kan du radera och skapa nya versioner.  
När du sparar en fil med versioner via kommandot Spara som... sparas inte versionsinformationen.  
Nya versioner  
Här skapar du nya versioner och / eller definierar om ytterligare en version ska skapas automatiskt när du stänger dokumentet.  
Spara ny version  
Om du klickar på den här kommandoknappen sparas dokumentet samtidigt som en ny version skapas.  
Innan du sparar kan du skriva en kommentar i en dialogruta.  
Mata in versionskommentar  
När du sparar en version skriver du in den kommentar du vill förse versionen med här.  
Du kan visa kommentaren till en sparad version genom att klicka på Visa men du kan inte redigera den.  
Spara alltid en version vid stängning  
Om den här rutan är markerad sparas alltid en version när dokumentet ändras och stängs.  
Då ställs alltid en kontrollfråga vid stängningen om det ändrade dokumentet ska sparas.  
Befintliga versioner  
Här listas alla befintliga versioner som du redan har skapat.  
Varje version förses med en tidsangivelse och innehåller information om författaren och en eventuell kommentar.  
Öppna  
Med den här kommandoknappen öppnar du den markerade versionen skrivskyddad i ett nytt fönster.  
Visa...  
Här kan du visa hela kommentaren till den markerade versionen.  
Radera  
Med denna markeras den valda versionen som raderad och dokumentet som modifierat.  
När du sparar dokumentet nästa gång raderas versionen verkligen.  
Jämför  
Med den här funktionen kan du jämföra de olika versionerna av dokumentet.  
Dialogrutan Acceptera eller ignorera ändringar öppnas.  
Ändringarna listas här och färgmarkeras i dokumentet.  
Ångra  
Med det här kommandot ångrar du den senaste åtgärden eller väljer åtgärden som du vill ångra i listrutan (som du öppnar genom att klicka längre med musen på ikonen).  
Bekräfta valet med returtangenten.  
För varje gång du klickar på ikonen upphävs den senaste åtgärden och så vidare.  
Antalet steg som du kan ångra ställer du in under Verktyg - Alternativ - %PRODUCTNAME - Arbetsminne.  
Observera att inte alla åtgärder (t.ex. ändringar av formatmallar) går att ångra med den här funktionen.  
Information för databastabeller  
För databastabeller är det bara möjligt att ångra den senaste åtgärden.  
Men detta gäller inte för databastabeller.  
När du redigerar databastabeller bör du tänka på följande: om du har ändrat innehållet i ett fält kan du ångra ändringen med ikonen Ångra.  
Om du ändrar fältinnehållet i en datapost som du ännu inte sparat, upphävs inte den senaste ändringen när ångra-funktionen används, utan processen "Inmatning av ny datapost", d.v.s. dataposten raderas i sin helhet.  
Information för presentationer  
När du väljer en ny sidlayout i en presentation måste listan med Ångra-åtgärder raderas.  
Ett meddelande informerar dig om detta och du kan eventuellt avbryta innan du väljer den nya sidlayouten.  
Återställ  
Med den här funktionen återställer du åtgärder som du tidigare har återkallat med Ångra.  
Om den senaste åtgärden inte ska återställas väljer du åtgärden som du vill återställa i listrutan (som du öppnar genom att klicka längre med musen på ikonen).  
Bekräfta valet med returtangenten.  
Senaste kommando  
Med denna funktion upprepas det sista kommandot.  
Du ser vilket kommando det är i menyn, efter menykommandot Senaste kommando.  
Klipp ut  
Med Klipp ut flyttar du det markerade objektet eller området till urklippet.  
Därifrån kan du infoga det i ett dokument hur många gånger du vill.  
Kopiera  
Det här kommandot kopierar det markerade objektet eller det markerade området till urklippet.  
Men om det redan finns ett innehåll i urklippet skrivs det över.  
Det går att använda urklippet med %PRODUCTNAME även i Unix-system.  
Men du måste använda %PRODUCTNAME -kommandona (Ctrl+C eller ikonen Kopiera på funktionslisten eller meny Redigera - Kopiera) när du vill kopiera från %PRODUCTNAME till urklippet.  
I det andra programmet räcker det sedan att trycka på musknappen i mitten.  
Om du vill kopiera från ett annat program räcker det att markera texten som skall kopieras och sedan välja kommandot i %PRODUCTNAME för att klistra in från urklippet (Ctrl+V eller ikonen Klistra in på funktionslisten eller meny Redigera - Klistra in).  
Klistra in  
Med detta kommando klistrar du in urklippets innehåll i dokumentet.  
I listrutan (som du öppnar genom att klicka längre på ikonen) kan du välja i vilket format innehållet i urklippet ska klistras in.  
Innehållet klistras in vid markörpositionen.  
Om en text eller ett objekt har markerats skrivs det markerade innehållet över av texten eller objektet som klistras in.  
Om ett område är markerat när celler kopieras från urklippet och om området är större än en rad resp. kolumn, men mindre än innehållet i urklippet, visas en dialogruta där du får en fråga om du verkligen vill utföra denna åtgärd.  
Om så är fallet klistrar programmet in utöver det markerade området.  
Klistra in innehåll Klistra in innehÃ¥ll  
Här bestämmer du i vilket format innehållet i urklippet ska klistras in i dokumentet.  
Urklippet kan innehålla olika datastrukturer, t.ex. text, bilder, grafik, tabellceller, ljudfiler m.m., men bara ett av dessa element åt gången.  
Via dialogrutan Klistra in innehåll kan du välja i vilket format innehållet i urklippet ska klistras in.  
Dialogrutan ser olika ut beroende på innehållet i urklippet.  
Om det finns celler från tabelldokument i urklippet visas en version av dialogrutan Klistra in innehåll, som beskrivs nedan.  
I alla andra fall visas den normala dialogrutan Klistra in innehåll som beskrivs först.  
Källa  
I det här visningsfältet ser du vilken typ av data som finns i urklippet, förutsatt att operativsystemet har kunnat definiera det.  
Urval  
I området Urval väljer du i vilket format som innehållet ska klistras in.  
Klistra in innehåll  
(Den här dialogrutan visas när data i urklippet kommer från tabellceller i tabelldokument.)  
Urval  
Det här området innehåller flera alternativ för vilket innehåll som ska infogas.  
Klistra in allt  
Om du markerar den här rutan klistras allt innehåll från det markerade cellområdet in.  
I annat fall skulle en senare ifyllning av de tomma cellerna i måldokumentet inte uppmärksammas.  
Strängar  
Om du markerar den här rutan infogas bara strängar.  
Siffror  
Om du markerar den här rutan infogas bara siffror.  
Datum och tid  
Om du markerar den här rutan infogas bara datum - och klockslagsposter.  
Formler  
Om du markerar den här rutan, infogas bara formler.  
Anteckningar  
Om du markerar den här rutan infogas bara anteckningar som du har lagt till i cellerna.  
Format  
Om du markerar den här rutan infogas bara de tilldelade formatattributen för celler.  
Räkneoperationer  
I det här området väljer du genom vilka räkneoperationer cellerna från urklippet ska kombineras med cellerna i det markerade målområdet.  
Den här funktion kräver att du markerar rutan Siffror i området Urval och ett område med celler i tabellen, där värden kan stå.  
De existerande värdena i målområdet kombineras med motsvarande värden från urklippet genom den valda räkneoperationen.  
Det är bara om en cell är tom i källområdet som behandlingen skiljer sig om du har valt funktionen Hoppa över tomma celler.  
Ingen  
Värdena från Urklipp infogas.  
Addera  
Värdena i Urklipp adderas till värdena i målområdet.  
Subtrahera  
Värdena i Urklipp subtraheras från värdena i målområdet.  
Multiplicera  
Värdena i urklippet multipliceras med värdena i målområdet.  
Dividera  
Värdena i målområdet divideras med värdena från Urklipp.  
Alternativ  
De här funktionerna reglerar på vilket sätt innehållet klistras in.  
Hoppa över tomma celler  
Om rutan Hoppa över tomma celler är markerad, påverkas inte den tillhörande målcellen när en tom rad "utan räkneoperation" infogas.  
Även när alternativet "Multiplicera" eller "Dividera "är markerat förändras inte målcellen.  
Om rutan Hoppa över tomma celler inte är markerad, tas alltså tomma rader med.  
En tom cell i källområdet raderar innehållet i motsvarande cell i målområdet om den infogas "utan räkneoperation".  
Vid multiplikation och division som räkneoperation behandlas en tom cell som en cell med innehåll 0.  
Det innebär att resultatet av multiplikationen alltid är 0 och resultatet av divisionen, om cellen i källområdet är tom, ger felmeddelandet #VÄRDE!.  
Transponera  
Om den här rutan är markerad transponeras innehållet i urklippet vid infogning; rader blir till kolumner och tvärtom.  
Länka  
Om du har markerat rutan Länka ändras det motsvarande värdet i målområdet när värdena i utgångsområdet ändras (som har kopierats till urklippet innan).  
Vill du också ta med senare ändringar av celler som för tillfället är tomma måste alternativet Klistra in allt vara markerat.  
Du kan också länka mellan tabeller i samma dokument.  
Om länkningen går utanför dokument skapas automatiskt en DDE-länk.  
En DDE-länk infogas som matrisformel och kan således bara ändras som helhet.  
Flytta celler  
Här definierar Du vad som ska hända med de existerande cellerna när det nya innehållet infogas.  
Flytta inte  
Markera det här alternativet när det infogade innehållet inte ska flytta de existerande cellerna.  
Nedåt  
Det här alternativet flyttar existerande celler i cellområdet nedåt när innehåll infogas.  
Höger  
Det här alternativet flyttar existerande celler i cellområdet åt höger när innehåll infogas.  
Markera allt  
Om du väljer menykommandot Markera allt markeras hela innehållet i den aktuella tabellen, det aktuella dokumentet, den aktuella ramen eller texten som har infogats som ritfunktion.  
Du kan också klicka på knappen utan text ovanför radhuvudena, till vänster om kolumnhuvudena.  
Du kan markera alla tabeller i ett dokument med kommandot Markera alla tabeller som finns på tabellflikarnas snabbmeny.  
Kommandon som används till en hel tabell gäller nu samtidigt för alla tabeller.  
Sök och ersätt  
Här kan du söka efter texter och / eller formateringar och ersätta dem med andra.  
Sök efter  
Här skriver du den text som du söker.  
Du kan öppna rutan och välja bland de senast angivna texterna.  
I området under Sök efter visas de valda attributen och formaten.  
Ersätt med  
Du kan öppna rutan och välja bland de senast angivna texterna.  
I området under Ersätt med visas de valda attributen och formaten.  
Alternativ  
Bara hela celler Bara hela ord  
Sökning sker efter celler vars innehåll exakt motsvarar sökordet.  
Om sökordet bara är en del av cellinnehållet hittas inte cellen.  
Om söktexten bara är en del av ett ord kommer den inte att hittas.  
Baklänges  
Sökningen börjar vid den aktuella markörpositionen och fortsätter mot dokumentets början.  
Reguljärt uttryck  
Markera Reguljärt uttryck om du vill använda platshållare i söktexten.  
Exakt sökning  
Om den här rutan är aktiverad måste texten stämma överens med söktexten när det gäller stor och liten bokstav för att den ska hittas.  
Bara markering  
Sökningen görs bara i texten som du har markerat.  
Sökning efter mallar  
Om den här rutan är markerad kan du söka efter celler som är formaterade med en viss cellformatmall.  
Vid Ersätt med kan du välja en ny cellformatmall som kan användas på de hittade cellerna.  
Välj styckeformatmallen vid Sök efter.  
Vid Ersätt med kan du välja en ny styckeformatmall som kan användas på de hittade styckena.  
Den här rutan heter Inklusive mallar när du har definierat ett attribut för sökningen med hjälp av knapparna Attribut eller Format.  
Markera den här rutan om du inte bara vill söka efter de direkta formateringarna utan även efter text som är formaterad med mallar som innehåller det attribut som du söker.  
Om du t.ex. söker efter attributet Språk så hittas normalt bara en effekt som du har använt direkt på tecken via Format - Tecken.  
Om du markerar rutan Inklusive mallar så hittas även de ställen där en teckenformatmall använts som bl.a. innehåller en definition av språket.  
Ta hänsyn till teckenbredd (bara om stödet för asiatiska språk är aktiverat)  
Om du klickar här tar sökningen hänsyn till halva / hela teckenbredder i asiatiska teckenuppsättningar.  
Likn. skrivsätt (japanska) (bara om stödet för asiatiska språk är aktiverat)  
Markera det här fältet om sökningen ska ta hänsyn till liknande skrivsätt på japanska.  
Via kommandoknappen... kommer du till en dialogruta där du kan göra de specifika inställningarna för likvärdig behandling och ignorering.  
Sök alla  
Startar sökningen.  
Alla träffar i hela dokumentet eller i markeringen som motsvarar söktexten och / eller attributen markeras.  
Sök  
Söker från och med den aktuella markörpositionen till nästa träff.  
Nästa träff är sedan markerad.  
Ersätt alla  
Alla träffar i dokumentet ersätts av ersättningstexten och / eller ersättningsattributen.  
När ersättningen är klar visas en dialogruta med antalet ersättningar som utförts.  
När du väljer kommandot Ersätt alla i %PRODUCTNAME Impress söks alla textblock igenom efter varandra, med början i det första textblocket.  
Om söktexten hittas i ett textblock ersätts den överallt i det här textblocket med ersättningstexten och sök-och-ersätt-operationen stoppas.  
Om du väljer kommandot på nytt söks nästa textblock igenom och så vidare till det sista textblocket.  
Till slut söks bakgrundssidorna igenom.  
När sökningen genom alla textblock och bakgrundssidor är avslutad meddelas det i en dialog.  
Ersätt  
Nästa träff ersätts av ersättningstexten och / eller ersättningsattributet.  
Attribut...  
Format...  
Inget format  
Klicka på den här kommandoknappen om du inte längre vill använda de valda attributen eller formaten för den fortsatta sökningen eller ersättningen.  
Klicka först i rutan vars attribut och format du vill stänga av (Sök efter eller Ersätt med) och klicka därefter på Inget format.  
De attribut som används visas under fälten.  
Fler>>  
Med den här kommandoknappen utökar du dialogrutan.  
Sök i  
Formler  
Det söks bara efter sökordet i formlerna.  
Du kan t.ex. hitta alla formler där SUMMA förekommer.  
Värden  
Det söks bara efter sökordet i värden.  
Du hittar t.ex. texter som bara beräknas och visas som resultat av en formel.  
Anteckningar  
Sökning sker endast i dokumentets anteckningar.  
Sökriktning  
Här väljer du mellan radvis eller kolumnvis sökriktning.  
Radvis  
Klicka här om du vill söka igenom tabellen radvis (horisontellt).  
Kolumnvis  
Klicka här om du vill söka igenom tabellen kolumnvis (vertikalt).  
Tillägg  
Sök i alla tabeller  
Markera den här rutan om du vill söka i alla tabeller i det aktuella dokumentet.  
Den här inställningen har högre prioritet än sökning bara i markerade tabeller.  
Fler<<  
Med den här kommandoknappen begränsar du dialogen.  
När du har stängt dialogrutan Sök och ersätt fortsätter du sökningen med hjälp av tangentkombinationen Skift Kommando +Ctrl +G.  
Du kan också fortsätta sökningen framåt och bakåt med hjälp av knapparna längst ned på den högra bildrullningslisten (vid den lilla Navigator-ikonen)  
Lista över reguljära uttryck  
Tecken  
Effekt / användning  
.  
Står för ett enda valfritt tecken.  
Om du skriver J.nsson hittar du "Jansson", "Jönsson" eller "Jonsson ".  
^Peter  
Ordet hittas enbart om det står i början av ett stycke.  
Särskilt innehåll (t.ex. tomma fält och ramar bundna till tecken) i början av ett stycke ignoreras.  
Peter$  
Ordet hittas enbart om det står i slutet av ett stycke.  
Särskilt innehåll (t.ex. tomma fält och ramar bundna till tecken) i slutet av ett stycke ignoreras.  
*  
Tecknet framför får förekomma hur många gånger som helst eller inte alls.  
Med Ab*c hittas t.ex. Ac, Abc, Abbc, Abbbc.  
För "valfria tecken eller inget tecken" kan man använda kombinationen .*  
+  
Tecknet framför måste förekomma minst en gång eller hur många gånger som helst.  
Med AX .+4 hittas AX 4, men inte AX4.  
Den längsta möjliga texten i ett stycke hittas alltid.  
Om texten AX 4 AX4 står i ett stycke, hittas den från det första A:et till den sista 4:an.  
?  
Med "Halv?" hittas orden "Hal "och "Halv".  
\C  
Exakt det här angivna tecknet (inga siffror) hittas, i det här fallet C (om du till exempel själv vill söka efter dollartecknet i ett reguljärt uttryck: \$)  
\n  
Hittar direkta radbrytningar som infogats med hjälp av Skift+Retur.  
Du kan också byta radbrytningar till styckebrytningar med hjälp av tecknet.  
Ange då \n både i fältet Sök efter och i fältet Ersätt med och bekräfta med kommandoknappen Ersätt alla.  
\t  
Hittar en tabb (det här uttrycket kan också stå i Ersätt med)  
\>  
Med "sol\>" hittas "vårsol "men inte "solsken".  
\<  
Med "\sol>" hittas "solsken "men inte "vårsol".  
^$  
Söker efter tomma stycken  
^.  
Söker efter första tecknet i ett stycke.  
&  
Med det här tecknet infogar du söktexten i fältet Ersätt med.  
Med "Fönster" i fältet Sök efter och "&båge "i fältet Ersätt med fås med hjälp av Ersätt "Fönsterbåge".  
Ange bara & i fältet Ersätt med om du vill tilldela söktexten andra Attribut eller ett annat Format.  
[abc123]  
Alla tecken som står inom parentesen hittas.  
[a-e]  
Alla tecken mellan a och e hittas  
[a-eh-x]  
Alla tecken i bokstavsgrupperna a-e och h-x hittas.  
[^a-s]  
Alla tecken utom a-s hittas  
\xXXXX  
Alla tecken med den fyrsiffriga hexadecimalkoden XXXX hittas  
Numret på ett tecken och även koden beror på det använda teckensnittet.  
Koderna finns under Infoga - Specialtecken.  
en _BAR_ ett  
Hittar alla "detta" och alla "det "  
{2}  
Det sista tecknet framför den inledande klammerparentesen måste förekomma så ofta efter varandra som siffran i parentesen anger.  
8{ 2} hittar 88.  
{1,2}  
Det sista tecknet framför den inledande klammerparentesen måste förekomma så ofta efter varandra som siffran i parentesen anger.  
8{ 1,2} hittar 8 och 88.  
()  
Med runda parenteser definierar du tecknen som står i parentesen som en referens.  
Sedan kan du använda den första referensen i det aktuella uttrycket med \1, den andra med \2 och så vidare.  
Om talet 13487889 står i din text och du söker efter det reguljära uttrycket (8 )7\1\1 hittas 8788.  
[:digit:]?  
Hittar en siffra (0 till 9).  
Med [:digit: ]* hittas en serie siffror.  
[:space:]?  
Hittar mellanrum som blanksteg och tabb.  
[:print:]?  
Hittar tecken som kan skrivas ut.  
[:cntrl:]?  
Hittar kontrolltecken.  
[:alnum:]?  
Hittar alfanumeriskt tecken (siffra och bokstav).  
[:alpha:]?  
Hittar alfabetiskt tecken (bokstav).  
[:lower:]?  
Hittar liten bokstav.  
[:upper:]?  
Hittar stor bokstav.  
Om du vill använda ett logiskt sökuttryck med kapslade OCH - / ELLER-operatorer använder du parenteser.  
Exempelvis söker du med "((a[A-z]*)_BAR_(ab[A-z]*)_BAR_(b[A-z]*))$" allt som börjar med ett mellanslag, fortsätter med "a "eller "ab" eller "b "och står i slutet av stycket.  
Likhetssökning  
Ställ in alternativen med hjälp av knappen....  
Den här sökningen skiljer sig från sökning med reguljära uttryck därför att den kan söka efter överensstämmelser på ett annat sätt.  
Den kan hitta ord som t.ex. skiljer sig åt från sökordet på två tecken som har bytt plats, infogats eller tagits bort på olika ställen.  
...  
Med den här kommandoknappen öppnas en dialogruta där du kan göra inställningar för likhetssökningen.  
Inställningar  
Här definierar du villkoren som ska gälla för att orden ska anses vara lika.  
Byt ut tecken  
Ange hur många tecken i sökordet som får vara utbytta för att en träff ska rapporteras.  
Vid standardinställningen på högst 2 tecken anses till exempel orden "skruv" och "strut "vara lika.  
Lägg till tecken  
Ange här hur många tecken längre ordet i dokumentet får vara jämfört med sökordet för att de fortfarande ska anses vara lika.  
Extratecknen får stå någonstans i ordet, i början, i slutet eller inne i ordet.  
Ta bort tecken  
Ange här hur många tecken kortare ordet i dokumentet får vara jämfört med sökordet, för att de fortfarande ska anses vara lika.  
Tecknen får tas bort från valfri plats i ordet, i början, i slutet eller inuti ordet.  
Kombinera  
Markera den här rutan om du vill kombinera de tre randvillkoren.  
Sökordet anses då vara funnet om ordet i dokumentet kan skapas genom en valfri kombination av de tre randvillkoren.  
Attribut  
Med den här kommandoknappen öppnar du en dialogruta där du kan välja attribut som ska sökas i den aktuella sökningen.  
Sökning sker efter alla direkta formateringar med attribut av den sökta typen, utan att du behöver specificera dem närmare.  
Om du väljer flera attribut så länkas de med ELLER.  
Om du vill söka efter särskilda attribut, exempelvis formatering med Courier, så klickar du på kommandoknappen Format  
Om du har definierat attribut ändras alternativrutan Sök efter formatmallar till Inklusive mallar.  
De aktuella, valda attributen räknas upp under textfältet Sök efter.  
Eftersom du kan välja fler attribut än vad som kan visas i det här fältet kan du placera markören i fältet och bläddra igenom de valda attributen med hjälp av piltangenterna.  
Om du inte bara vill söka efter direkta formateringar utan även formateringar som har gjorts med formatmallar med de här attributen markerar du rutan Inklusive mallar i området Alternativ.  
Urval  
Här väljer du de attribut som du vill söka efter.  
Håll ihop stycken  
Här söker du efter attributet Håll ihop stycken.  
Dela stycke  
Här söker du efter attributet Dela inte stycke.  
Avstånd  
Här söker du efter attributet Avstånd (Uppe, Nere).  
Justering  
Här söker du efter attributet Justering (Vänster, Höger, Centrerat, Marginaljustering).  
Effekter  
Här söker du efter effekterna Små kapitäler, Versaler, Titelteckensnitt och Gemener.  
Blinkande  
Här söker du efter attributet Blinkande.  
Genomstruken  
Här söker du efter attributet Genomstruken (enkelt eller dubbelt).  
Indrag  
Här söker du efter attributet Indrag (Från vänster, Från höger, Första raden).  
Horungar  
Här söker du efter attributet Horungekontroll.  
Kerning  
Här söker du efter attributen Avstånd (Standard, Spärrat, Smalt) och parvis Kerning.  
Kontur  
Här söker du efter attributet Kontur.  
Position  
Här söker du efter positionen Normal, Upphöjd eller Nedsänkt.  
Register  
Här söker du efter attributet Register.  
Relief  
Här söker du efter attributet Relief.  
Rotation  
Här söker du efter attributet Rotation.  
Skuggad  
Här söker du efter attributet Skugga.  
Teckensnitt  
Här söker du efter attributet Teckensnitt (teckensnittets namn).  
Teckenfärg  
Här söker du efter en teckenfärg.  
Teckenstorlek  
Här söker du efter attributet Teckenstorlek / teckenhöjd.  
Tjocklek  
Här söker du efter attributet Fet eller Fet Kursiv.  
Teckenstil  
Här söker du efter attributet Kursiv eller Fet Kursiv.  
Änkor  
Här söker du efter attributet Änkekontroll.  
Sidformatmall  
Här söker du efter attributet Brytning med sidformatmall.  
Avstavning  
Här söker du efter attributet Avstavning.  
Skalning  
Här söker du efter attributet Skalning.  
Språk  
Här söker du efter attributet Språk (för rättstavningskontroll).  
Tabulatorer  
Här söker du efter ett stycke som innehåller en extra tabb.  
Understruken  
Här söker du efter attributet Understruken (enkelt, dubbelt eller punkterat).  
Vertikal textjustering  
Här söker du efter attributet Vertikal textjustering.  
Ordvis  
Här söker du efter attributet Ordvis (när det är understruket eller genomstruket).  
Teckenbakgrund  
Här söker du efter attributet Teckenbakgrund.  
Radavstånd  
Här söker du efter attributet Radavstånd (Enkelt, 1,5 rad, Dubbelt, Proportionellt, Minst, Eget radavstånd).  
Textattribut  
Detta skiljer sig från sökningen med hjälp av kommandoknappen Attribut... då du söker efter alla attribut av den valda typen.  
De aktuella, valda attributen räknas upp under textfältet Sök efter.  
Eftersom Du kan välja fler attribut än vad som kan visas i detta fält kan Du placera markören i fältet och bläddra igenom de valda attributen med hjälp av piltangenterna.  
Om du bara vill söka och ersätta särskilda attribut, oberoende av texten, raderar du det om står i textfältet Sök efter.  
Du definierar attributen för ersättningen genom att först klicka i textfältet Ersätt med och därefter välja Format.  
I båda fallen definierar du attributen i dialogrutan Textattribut.  
I den här dialogrutan finns följande flikar.  
Navigator för samlingsdokument  
När du har öppnat ett samlingsdokument kan du växla mellan normalläge och samlingsläge för Navigator.  
I visningsfältet listas alla poster i samlingsdokumentet.  
Här kan Du även kontrollera om det finns länkar till alla de deldokument som visas.  
Håll muspekaren över en valfri post så visas sökvägen till det länkade dokumentet.  
Om t ex ett originaldokument har tagits bort, dvs inte finns kvar på den ursprungliga platsen, visas meddelandet Hittar inte filen i rött tillsammans med sökvägen.  
I samlingsläget visas inte listrutan Öppnade dokument i Navigator och antalet och typ av ikoner varierar:  
Växla  
Med den här ikonen växlar du mellan samlingsläge och normalläge för Navigator.  
Växla  
Redigera  
Markera en post i Navigator och klicka här för att redigera innehållet.  
Om den markerade posten är en fil öppnas det länkade dokumentet för redigering, är den en förteckning öppnas en dialogruta för förteckningar, är den en text placeras markören i textstycket.  
Redigera  
Uppdatera  
Här öppnas en undermeny där du väljer vilket innehåll som ska uppdateras.  
Du kan välja det markerade innehållet, befintliga förteckningar, alla länkar eller samtliga poster.  
Uppdatera  
Markering  
Det markerade innehållet uppdateras.  
Förteckningar  
Förteckningarna uppdateras.  
Länkar  
Länkarna uppdateras.  
Allt  
Allt innehåll uppdateras.  
Redigera länk  
Det här kommandot på en snabbmeny i ett infogat dokument öppnar dialogrutan Redigera områden Redigera områden.  
Infoga  
Klicka här om du vill infoga en förteckning, ett dokument eller en text i samlingsdokumentet.  
Då öppnas en undermeny med aktuella alternativ.  
Du kan också infoga filer i samlingsdokumentet genom att dra och släppa dem med musen.  
Sedan öppnas det och du kan redigera och spara det direkt.  
Infoga  
Förteckning  
Med det här kommandot kan Du infoga en valfri förteckning.  
Fil  
Med det här kommandot öppnar Du en dialogruta i vilken Du kan infoga en fil.  
Nytt dokument  
Med det här kommandot skapar Du ett nytt textdokument.  
Först visas dialogrutan Spara som där Du kan ge det nya dokumentet ett namn och bestämma var det ska sparas.  
Text  
Med det här alternativet placerar Du markören i samlingsdokumentet, och Du kan därefter skriva in text.  
Spara med innehåll  
När den här knappen är intryckt sparas innehållet i de länkade filerna även i samlingsdokumentet.  
Det tar dubbelt så stor plats, men innehållet är då tillgängligt även om de länkade filerna inte är det.  
Spara med innehåll  
Flytta nedåt  
Klicka på den här ikonen om du vill flytta den markerade posten nedåt i Navigator-rutan.  
Du kan även flytta poster med dra-och-släpp.  
Om textområden flyttas ihop sammanfogas de till ett enda textområde.  
Flytta nedåt  
Flytta uppåt  
Klicka på den här ikonen om du vill flytta den markerade posten uppåt i Navigator-rutan.  
Du kan också flytta poster genom att dra och släppa dem.  
Om textområden flyttas ihop sammanförs de till ett enda textområde.  
Flytta uppåt  
Radera  
Med det här kommandot raderar du den markerade posten i visningsfältet i Navigator.  
Redigera länkar  
Här kan du redigera de länkar som fogats in i det aktuella dokumentet.  
Den här funktionen kan bara användas om det aktuella dokumentet innehåller länkar.  
I dialogrutans listruta listas de länkar som finns i det aktuella dokumentet.  
Information om sökväg och filnamn för en länk bibehålls även om den länkade datafilen inte finns på den använda datorn, eller om den flyttas till en annan katalog.  
Så snart den länkade filen finns tillhands på det angivna stället kan den också användas i dokumentet.  
När du öppnar en fil som innehåller länkar får du en fråga om länkarna ska uppdateras nu.  
På så sätt betraktas inga länkar av misstag som kontrollerade under genomgången, som kan ta ganska lång tid med långsamma servrar.  
Vid laddningen av filer som innehåller DDE-länkar får Du en fråga om länken ska uppdateras.  
Du kan svara Nej på detta om Du inte vill att DDE-servern ska anropas.  
Källfil  
Här visas den länkade filens URL.  
Element  
Här visas den länkade filens typ och eventuellt också det program med vilken filen skapades.  
Typ  
Den länkade filens typ (grafik, text osv) visas här.  
Status  
Under listrutan visas information om den markerade länken.  
Automatisk  
Om den länkade datafilen uppdateras genomför programmet den nödvändiga uppdateringen.  
Denna uppdateringsmetod är meningsfull om Du hela tiden vill arbeta med den länkade datafilens senaste version.  
Vid länkade grafikobjekt är detta fält inte aktivt, eftersom grafikobjekt bara kan uppdateras manuellt.  
Manuellt  
Uppdateringen måste utföras av användaren.  
Denna uppdateringsmetod är meningsfull om Du själv vill bestämma när Du vill använda den senaste versionen av den uppdaterade filen i Ditt dokument.  
Vid länkade grafikobjekt är detta fält inte aktivt, eftersom grafikobjekt bara kan uppdateras manuellt.  
Uppdatera  
Den eller de markerade filernas länkar uppdateras.  
Nu visas den senaste versionen av den eller de länkade filerna.  
Efter uppdateringen visas återigen den första markerade posten.  
Ändra  
Om Du vill ersätta den aktuella länkade filen med en annan fil eller ändra sökvägen till länkningen använder Du denna kommandoknapp.  
Sökvägen respektive filen ändras med en standarddialog för val av filer (med undantag för DDE-länkar).  
Vid en befintlig DDE-länk kommer Du till dialogrutan Ändra länk.  
Upplös  
Hänvisningen till filen tas bort ur dokumentet.  
Denna åtgärd är meningsfull om Du bara vill arbeta med den senaste versionen av den länkade filen, eller om dokumentet ska redigeras på en annan dator och den länkade filen inte kan kopieras till den andra datorn.  
Innan länkens upplöses får Du en kontrollfråga.  
Ändra länk  
I den här dialogrutan visas de aktuella parametrarna för den markerade DDE-länken och du kan ändra dem.  
Ändra länk  
I det här området visas de parametrar som för tillfället gäller för länken.  
Applikation:  
I det här fältet kan Du växla program, om DDE-länken hänför sig till ett annat program.  
Fil:  
Här visas länkens aktuella sökväg.  
Område:  
Om du vill byta det område som länken ska hänvisa till, skriver Du in det här.  
Plug-in  
Med det här kommandot aktiverar eller deaktiverar du plug-ins (insticksprogram).  
Om en plug-in är aktiv kan den inte flyttas i dokumentet eller redigeras utan måste deaktiveras först.  
Objekt  
Med det här kommandot kan du redigera ett infogat objekt.  
Du kan bara använda det här kommandot om minst ett objekt är infogat i dokumentet. (Se Infoga - Objekt)  
Om du vill redigera eller öppna ett objekt som är infogat i dokumentet, måste du först markera det genom att klicka på det.  
En undermeny öppnas som innehåller följande funktioner:  
Redigera  
Med det här kommandot kan du redigera ett infogat objekt.  
Om du vill redigera ett objekt, markerar du det först och väljer sedan det här kommandot.  
Då visas verktygen med vilka du kan redigera det markerade objektet.  
Detta fungerar bara med %PRODUCTNAME -objekt.  
Om du t.ex. vill redigera ett MS-Excel-objekt, måste du använda Excel.  
Om ett objekt infogas via OLE, så är det objektet som registrerar denna menypost i %PRODUCTNAME -programmets meny.  
Öppna  
Med det här kommandot öppnas objektet med det program med vilket det ursprungligen skapades.  
Där kan du redigera det.  
Objektet visas i ett separat dokumentfönster.  
Detta menykommando infogas i menylisten av det program som är länkat till objektet som ska redigeras.  
Därför kan kommandot även heta något annat, t ex Open.  
Nedanför objektlisten visas redigeringsprogrammets funktionslist.  
När alla ändringar är gjorda stänger Du dokumentfönstret med ikonen Stäng på titellisten.  
Det inbäddade objektet uppdateras.  
Om Du vill kunna använda denna funktion måste Du ha infogat objektet via menyn Infoga och kommandot Objekt.  
Ram - egenskaper  
I den här dialogrutan anger du grundläggande egenskaper för en ram.  
Namn  
I det här textfältet ger du ramen ett namn.  
Namnet måste uppfylla kraven för namn i HTML-språket och bör alltså bara bestå av tecknen a till z och 1 till 0 (inte å, ä, ö, inga blanksteg).  
Namn med understreck (_) i början är reserverade namn som du inte får använda själv.  
Innehåll  
I det här textfältet anger du URL:n för filen som du vill lägga till i den aktuella ramen.  
Exempel:  
http: / /www.sun.se  
file: / //c _BAR_ / Laesmig.txt  
Du kan också använda... till höger om textfältet och söka efter URL:n.  
...  
Om du klickar på den här kommandoknappen, öppnas dialogrutan Välj ut fil för ram.  
Den motsvaras av dialogrutan Arkiv - Öppna.  
Välj filen som du vill lägga till i den aktuella ramen.  
Rullningslist  
I det här området bestämmer du om den aktuella ramen ska ha en vertikal rullningslist.  
På  
Välj det här alternativet om ramen alltid ska ha en rullningslist.  
Av  
Välj det här alternativet om den aktuella ramen aldrig ska ha en rullningslist.  
Du måste då rulla genom innehållet med piltangenterna om det inte passar in i ramen.  
Automatiskt  
Välj det här alternativet om den aktuella ramen ska få en rullningslist vid behov.  
Inramning  
Här väljer du typ av inramning.  
På  
Välj det här alternativet om ramen ska ha en synlig kant.  
Av  
Välj det här alternativet om ramen inte ska ha någon synlig kant.  
Avstånd till innehåll  
I det här området anger du hur mycket plats som ska finnas mellan kanten på en ram och ramens innehåll, eller så använder du standardinställningarna.  
Bredd  
Här definierar du det horisontella avståndet mellan ramens innehåll och kant.  
Höjd  
Här definierar du det vertikala avståndet mellan ramens innehåll och kant.  
Standard  
Om du markerar den här rutan används standardinställningarna för respektive avstånd.  
Image map-redigerare  
Med den här redigeraren kan du skapa klickbara grafikobjekt.  
Definiera de områden inom ramar och grafikobjekt som ska utlösa speciella åtgärder när man klickar på dem.  
Till varje område inom ramen eller grafikobjektet kan Du koppla en URL, som ska laddas när Du klickar på detta område i ImageMap en.  
Du anger om den nyladdade URL:en ska visas i ett eget fönster, i samma fönster eller i en ram.  
På de överlappande ställena gäller det sist definierade området.  
Vid målen kan du välja helt fritt om de t.ex. ska hänvisa till Internet-sidor eller referenser i det aktuella dokumentet eller i ett annat dokument i filsystemet.  
Tilldela  
Efter varje ny post och efter varje ändring av en post i image map-redigeraren klickar du på den här ikonen för att tilldela den aktuella ändringen.  
Tilldela  
Öppna  
Klicka här om du vill öppna en image map-fil i filformaten MAP-CERN, MAP-NCSA eller SIP StarView ImageMap.  
Öppna  
Spara  
Sparar image map i något av filformaten MAP-CERN, MAP-NCSA eller SIP StarView ImageMap.  
En dialogruta visas där du kan spara en fil.  
Spara  
Urval  
Klicka på ikonen Urval så aktiveras urvalsmarkören.  
Med den här markören kan du markera en annan del i en image map för att sedan redigera den.  
Urval  
Rektangel  
Klicka på Rektangel om du vill definiera ett rektangulärt område.  
Markören får en liten rektangel bredvid hårkorset och du kan nu rita upp en rektangel med musen.  
Om du vill skapa en kvadrat håller du ner skifttangenten samtidigt som du drar.  
När du släpper musknappen kan du mata in uppgifter för det här området i fälten Adress, Text och Frame.  
Rektangel  
Ellips  
Klicka på Ellips om du vill definiera ett runt område.  
Markören får en liten cirkel bredvid hårkorset och du kan nu rita upp en ellips med musen.  
Om du vill skapa en cirkel håller du ner skifttangenten samtidigt som du drar.  
När du släpper musknappen kan du mata in uppgifter för det här området i fälten Adress, Text och Frame.  
Ellips  
Polygon  
Klicka på Polygon om du vill definiera ett fritt område.  
Markören får en liten kurva bredvid hårkorset och du kan nu definiera en polygon.  
Klicka på varje punkt på kurvan som du vill definiera.  
Dubbelklicka på startpunkten för att sluta kurvan.  
Du kan begränsa vinkeln till multiplar av 45 grader om du håller ner skifttangenten när du placerar muspekaren.  
När du har slutit kurvan kan du mata in uppgifter för området i fälten Adress, Text och Frame.  
Polygon  
Frihandspolygon  
Klicka på Frihandspolygon om Du vill definiera ett valfritt område.  
Markören får en liten kurva bredvid hårkorset och Du kan nu definiera en frihandspolygon.  
Klicka på kurvans startpunkt och dra med nedtryckt musknapp ut det område som Du vill definiera.  
När Du släpper musknappen sluter sig polygonen automatiskt.  
Frihandspolygon  
Redigera punkter  
Klicka på Redigera punkter om Du vill visa enstaka stödpunkter på Bézierkurvor.  
Då kan Du redigera de enskilda stödpunkterna på kurvan med hjälp av musen.  
Redigera punkter  
Flytta punkter  
Klicka på Flytta punkter om Du vill flytta enstaka punkter som definierar en polygon.  
Flytta punkter  
Infoga punkter  
Klicka på Infoga punkter om Du vill infoga ytterligare stödpunkter.  
Infoga punkter  
Ta bort punkter  
Klicka på Ta bort punkter om Du vill ta bort enstaka stödpunkter.  
Ta bort punkter  
Aktiv  
Med den här ikonen växlar du mellan aktivt och inaktivt läge för den markerade delen av image map.  
Den här funktionen behöver du normalt inte använda när du skapar en image map utan först senare när du ska uppdatera ett sådant grafiskt objekt.  
Då behöver Du inte skapa hela det grafiska objektet på nytt.  
En inaktiv ram är i motsats till en aktiv transparent.  
Aktiv  
Makro  
När du klickar på den här ikonen visas dialogrutan Tilldela makro, som är uppbyggd på samma sätt som dialogrutan Makro.  
Här tilldelar du en image map ett makro.  
Makro  
Egenskaper  
Om du klickat på den här ikonen öppnas dialogrutan Beskrivning, där du kan definiera URL, Alternativtext, Ram och Namn.  
Egenskaper  
Adress:  
Markera i detta kombinationsfält den URL (eller lokala fil) som ska laddas då Du klickar på området.  
Referenser inom filen läggs till filnamnet enligt skrivsättet för URL.  
Om Du t ex vill hoppa till ankaret "Här" (som Du har definierat med Infoga - Fältkommando - Andra - Referenser - Sätt referens) i filen C:\Docs\Test.sdw anger Du adressen: file: / //C _BAR_ / Docs / Test.sdw#Här.  
Text:  
Den text Du anger här visas när Du pekar med musen på området i grafiken.  
Om det inte finns någon text visas adressen.  
Denna text motsvarar fältet Alternativtext i dialogrutan Beskrivning.  
Ram:  
Här markerar Du den målram som det anropade dokumentet ska laddas i.  
Förklaringstabell  
Grafikvy  
Här kan du definiera konturerna som ska reagera på ett visst sätt när man klickar på dem.  
Beskrivning  
I den här dialogrutan finns information om URL, alternativtext, ramtyp och namnet på det markerade området i grafiken.  
Hyperlänk  
Här finns all information om hyperlänken.  
URL:  
I det här textfältet anger Du den URL (eller lokala fil) som ska laddas då Du klickar på området.  
Referenser inom filen läggs till filnamnet enligt skrivsättet för URL.  
Om Du till exempel vill hoppa till ankaret "Här" (som Du har definierat med Infoga - Fältkommando - Andra... - Referenser - Ställa in referens) i filen C:\Docs\Test.sdw, anger Du följande adress: file: / //C _BAR_ / Docs / Test.sdw#Här.  
Alternativtext:  
Den text du anger här visas när du pekar med musen på grafikområdet.  
Om det inte finns någon text visas adressen.  
Detta fält motsvarar fältet Text i Image map-redigeraren.  
Ram:  
Här markerar du ramen som dokumentet ska laddas i.  
De förinställda posternas betydelse hittar du i förklaringstabellen.  
Namn:  
Här tilldelar Du det markerade området i grafiken ett namn.  
Ändringar  
Här hittar du olika kommandon för registrering och visning av ändringar i dokument.  
Du kan skriva kommentarer till registrerade ändringar.  
Visa  
Visa  
Acceptera eller ignorera...  
Kommentar...  
Sammanfoga dokument...  
Registrera  
Med det här kommandot startar eller avslutar du registreringen av en ändring i ett dokument.  
Om du har aktiverat funktionen Registrera finns en bock framför menykommandot.  
Ändringar som du gör i dokumentet registreras från och med nu tills du avslutar registreringen genom att åter aktivera kommandot.  
De ställen som du har ändrat markeras med ett streck i marginalen om du har markerat både Registrera och Visa.  
Egenskaperna för strecket ställer du in under Verktyg - Alternativ - Textdokument - Ändringar.  
Registreringen omfattar följande ändringar av dokumentinnehållet:  
Infoga och radera text  
Flytta stycken  
Sortera text  
Söka och ersätta text  
Infoga attribut som är ett tecken brett, t.ex. fält och fotnoter  
Infoga tabeller, områden  
Infoga dokument  
Infoga AutoText  
Infoga via urklipp  
Ändra cellinnehåll med hjälp av infogning och radering  
Infoga eller radera kolumner och rader  
Infoga tabellark  
Klippa ut, kopiera och infoga via urklippet  
Flytta med dra-och-släpp  
Ändringar i formler eller tal i tabeller registreras inte.  
Medan registreringen är aktiverad kan du inte radera, flytta eller kopiera tabeller.  
De enskilda ändringarna behandlas som infogningar respektive raderingar och förs in i en ändringslista.  
Du styr visningen av de registrerade ändringarna i dokumentet med menykommandot Visa.  
Du anger hur ändringarna i dokumentet ska visas under Verktyg - Alternativ - Textdokument... - Ändringar.  
Du anger hur ändringarna i dokumentet ska visas under Verktyg - Alternativ - Tabelldokument... - Ändringar.  
Skydda registrering  
Här skyddar du registrerade ändringar genom att ange ett lösenord.  
Samtidigt aktiveras registreringen av ändringar.  
Om Skydda registrering är aktiverat går det bara att stänga av registreringen igen med det här kommandot och det riktiga lösenordet.  
Visa ändringar  
Här anger du om registrerade ändringar i dokumentet ska visas.  
Om du har aktiverat funktionen Visa finns det en bock framför menykommandot.  
Alla ändringar har som registrerats eller som du just registrerar visas då i dokumentet.  
Registrerade ändringar framhävs i färg i tabellen.  
Under Verktyg - Alternativ - Tabelldokument... - Ändringar definierar du färgerna för de olika ändringarna.  
I standardinställningen är inmatningar understrukna och raderingar genomstrukna.  
Du kan ändra dessa inställningar under Verktyg - Alternativ - Textdokument... - Ändringar.  
En ändring sparas alltid tillsammans med följande information: uppgifter om författaren som har gjort ändringarna hämtas från de användardata som finns i %PRODUCTNAME (Verktyg - Alternativ - %PRODUCTNAME - Användardata).  
Datum och klockslag för ändringen hämtas från systeminställningarna.  
Du kan ange en kommentar till ändringen under Redigera - Ändringar - Kommentar.  
Författare, datum och klockslag för ändringen visas i tips-hjälpen när du för musen över den markerade ändringen i dokumentet.  
Om du har slagit på den aktiva hjälpen visas dessutom kommentaren.  
Vidare visas ändringens typ och innehåll.  
Visa ändringar i tabellen  
Markera det här fältet när ändringar i tabellen ska visas.  
Visa accepterade ändringar  
Tillhörande kommentarer visas också.  
Visa ej accepterade ändringar  
Tillhörande kommentarer visas också.  
Kommentera ändring  
Du kan titta på en befintlig kommentar och vid behov redigera den.  
Du kan också använda funktionen när du har markerat en ändring om du öppnar snabbmenyn i dialogrutan Acceptera eller ignorera ändringar och väljer Redigera kommentar... Redigera kommentar  
Kommentarer visas precis som för anteckningar i en förklaring i tabelldokumentet samt i ändringslistan i dialogrutan Acceptera eller ignorera ändringar.  
Dialogrutan där du kan skriva eller redigera en kommentar motsvarar dialogrutan för Infoga anteckning.  
Acceptera eller ignorera ändringar  
Här visas dialogrutan där du accepterar eller avböjer enskilda ändringar i ett dokument.  
Lista  
Där finns också ytterligare information.  
På denna sida På denna flik finns en förteckning över alla ändringar som uppfyller de inställda filterkriterierna.  
Det finns dock ett undantag.  
Då ändringarna är kapslade visas beroenden oberoende av vilket filter som har angetts.  
Kapslade ändringar är sådana där olika åtgärder för ett textställe delvis sammanfaller.  
Det kan t ex vara när flera författare gör ändringar på samma ställe i texten.  
Antag att författare A infogar en text i ett dokument och att författare B raderar en del av denna text.  
Detta beror på att den ursprungliga infogningen från författare A inte längre motsvarar det aktuella dokumentet.  
Om flera ändringar har gjorts i samma cell visas alla dessa ändringar som en enda post i listan.  
Klicka på plustecknet bredvid posten om Du vill se mer detaljerade uppgifter om de enskilda ändringarna.  
Om flera ändringar ha gjorts i en cell kommer alla ändringar att visas, oberoende av vilka filterkriterier som Du har ställt in, om åtminstone en av ändringarna uppfyller filterkriterierna.  
De olika posterna i ändringslistan är färgmarkerade om Du har angett ett filter.  
De olika färgerna har följande betydelser:  
Färg  
Betydelse  
svart  
Posten kan accepteras, avböjas och motsvarar filterkriterierna.  
blå  
Posten kan accepteras, avböjas men motsvarar själv inte filterkriteriet.  
Det finns dock en eller flera underposter som motsvarar kriteriet.  
grå  
Underposten kan inte accepteras eller avböjas samt motsvarar inte filterkriteriet.  
grön  
Underposten kan inte accepteras eller avböjas men motsvarar filterkriteriet.  
Listruta  
Här visas ändringarna.  
När du markerar en post i listan visas motsvarande ändring i dokumentet.  
Du kan också markera flera poster samtidigt med hjälp av Ctrl-tangenten.  
Du kan också acceptera resp. avböja alla ändringar på en gång.  
Du kan t ex sortera listan genom att klicka på kolumnrubrikerna, ställa in optimal bredd genom att dubbelklicka på skiljelinjen mellan kolumnrubrikerna osv.  
I en posts snabbmeny finns ytterligare kommandon för att ändra sorteringen och redigera kommentarer.  
När du har accepterat eller avböjt en ändring sorteras listposterna hierarkiskt efter "Accepterade" och "Tillbakavisade ".  
Åtgärd  
Här visas i klartext vilken åtgärd som beskrivs i den här posten.  
Position  
Här visas vilken eller vilka celler respektive områden som berörs av ändringen.  
Författare  
Här visas vem som har gjort ändringen.  
Datum  
Här visas datumet för ändringen.  
Beskrivning  
Här visas en exakt beskrivning av ändringen.  
Acceptera  
Klicka här om du vill acceptera den markerade posten.  
Avböj  
Klicka här om du vill avböja den markerade posten.  
Ändringen ignoreras då slutgiltigt och det ursprungliga innehållet återställs.  
Acceptera alla  
Klicka här om du vill acceptera alla ändringar.  
Avböj alla  
Klicka här om du vill avböja alla ändringar.  
Ändringar som du har accepterat eller avböjt kan tas tillbaka med menykommandot Redigera - Ångra.  
Ångra  
Om du har skapat och registrerat ändringar med hjälp av AutoFormat-funktionen (menykommandot Format - AutoFormat - Använd och redigera ändringar)), innehåller dialogrutan dessutom kommandoknappen Ångra.  
Alla ändringar som du har gjort med AutoFormat listas en och en och du kan acceptera respektive ignorera varje enskild ändring.  
Med hjälp av kommandoknappen Ångra kan du återställa ändringar som du har accepterat eller ignorerat.  
Det finns fler kommandon på listans snabbmeny:  
Redigera kommentar  
Här kan du skriva och redigera en kommentar (som visas i kolumnen Beskrivning).  
Sortera efter  
En undermeny öppnas där du kan välja vilken kolumn som listan ska sorteras efter.  
Åtgärd  
Listan sorteras efter typ av åtgärd.  
Författare  
Listan sorteras efter författare.  
Datum  
Listan sorteras efter datum.  
Beskrivning  
Listan sorteras efter kommentar.  
Dokumentposition  
Listan sorteras, uppifrån och ned, efter ändringens position i dokumentet Detta är standardinställningen.  
Filter  
Här anger du vilka ändringar du vill se - av vilken författare och från vilken tidsperiod.  
De filtervillkor som ställts in under den här fliken avgör vilka ändringar som ska föras in under fliken Lista.  
Datum  
Ange tidsperioden i fälten nedanför.  
Om rutan inte är markerad, kommer alla ändringar som hittills är gjorda att visas.  
Ställ in datum / klockslag  
Om du klickar på den här ikonen anges automatiskt aktuellt datum och klockslag i respektive fält.  
Författare  
Om bara ändringarna som har gjorts av en viss person ska visas, markerar du den här rutan och väljer i kombinationsfältet den författare vars ändringar du vill se.  
Om rutan inte är markerad, kommer alla ändringar att visas oavsett vem som har gjort dem.  
Område  
Ange området i textfältet.  
Du kan också använda funktionen Ställ in tabellreferens när du ska ange området.  
Om rutan inte är markerad, visas alla ändringar i hela tabelldokumentet.  
Ställ in tabellreferens  
Om du klickar på den här kommandoknappen, kan du markera önskat tabellområde med musen.  
Tabellreferensen förs då in i textfältet.  
Om du klickar på kommandoknappen, minimeras dialogrutan.  
Markera det tabellområde vars ändringar du vill se och förstora sedan dialogrutan genom att klicka på motsvarande ikon.  
Förminska / Förstora  
När du har markerat ett område i tabellen med musen, klickar du på den här ikonen om du vill återställa dialogrutan till ursprunglig storlek.  
Åtgärd  
Välj sedan önskad åtgärd i kombinationsfältet.  
Om rutan inte är markerad, visas alla åtgärder.  
Beskrivning  
Du kan filtrera visningen av ändringar enligt särskilda beskrivningar.  
De beskrivningarna visas i listan över ändringar.  
Du får information om typen av ändring och eventuell tillhörande kommentar.  
Markera kryssrutan Beskrivning om bara de ändringar ska visas vars beskrivning innehåller en viss text, som Du anger i textfältet intill.  
Om Du t ex vill se alla ändringar som i kommentaren innehåller ordet "viktigt", skriver Du "viktigt" under Beskrivning.  
När Du ska filtrera enligt särskilda beskrivningar kan Du också använda platshållare.  
Du kan därvid använda samma reguljära uttryck som i dialogrutan Sök och ersätt.  
Infoga (Sammanfoga dokument)  
Då kan Du i det aktuella dokumentet (originaldokumentet) klistra in de ändringar som har gjorts i en kopia av det dokumentet.  
I det aktuella dokumentet visas då de textställen det cellinnehåll som är identiskt lika i det aktuella och det inklistrade dokumentet i bara en uppsättning, medan varje del som har ändringsmarkerats i något av dokumenten visas.  
Förutom innehållet hämtas också uppgifter om ändringarnas författare och datum samt tillhörande kommentarer.  
Förutsättningen för att det gå att sammanfoga två dokument är att båda har samma ursprung, d.v.s. de får bara skilja sig åt i fråga om ändringarna.  
På det här sättet kan du sammanfoga flera kopior av ett dokument till ett enda dokument alltefter behov.  
För närvarande är det bara den löpande texten som sammanfogas, dvs inte fotnoter, sidhuvuden eller sidfötter, ramar eller fält.  
Infoga (Jämför dokument)  
Välj ett dokument som ska jämföras med det aktuella dokumentet.  
Skillnaderna mellan dokumenten markeras som ändringar i det aktuella dokumentet.  
För närvarande jämförs bara den löpande texten, d.v.s. inte fotnoter, sidhuvuden eller sidfötter, ramar eller fält.  
Litteraturdatabas  
Med det här kommandot kan du infoga nya dataposter i litteraturdatabasen och redigera befintliga data.  
Litteraturdatabasen innehåller ett antal dataposter med information om böcker om %PRODUCTNAME.  
I en gemensam vy med dataposterna i tabellform och markerade dataposter i ett formulär.  
Med hjälp av objektlisten kan du välja en viss tabell i bibliografidatabasen, söka efter innehåll och använda filter.  
Välja ut datapost  
Välja ut tabell  
Välj ut tabellen som innehåller den sökta dataposten i listrutan.  
Gå till datapost  
Det finns flera kommandoknappar som Du använder när Du vill gå till en datapost i tabellen  
Hopp till den första dataposten i tabellen.  
Hopp till föregående datapost.  
Hopp till nästa datapost.  
Hopp till den sista dataposten i tabellen.  
Om Du vet numret på den sökta dataposten kan Du mata in det i datapostfältet för att komma till dataposten.  
Infoga ny datapost  
Klicka på den här kommandoknappen om Du vill skapa en ny datapost.  
Klicka på ikonen med en asterisk (*) på datapostlisten (i tabellvyns undre kant).  
En ny, tom rad skapas och visas i tabellen, och inmatningsmarkören placeras i det första datafältet.  
Klicka i listrutan Typ i formuläret som finns i nedre delen av fönstret.  
Välj typ av litteraturhänvisning.  
I det första fältet anger Du den korta beteckningen som ska stå som referens i Ditt textdokument.  
Mata in de andra uppgifterna för den nya dataposten i formuläret.  
Innehållet i ett datafält sparas automatiskt när du flyttar markören till ett annat datafält i samma datapost.  
Filtrera och söka dataposter  
Textfältet Sökbegrepp och filterikonerna används till att söka innehåll i tabellen.  
Mata in sökbegrepp  
Mata in ett sökbegrepp i textfältet.  
Alla dataposter som börjar exakt likadant som sökbegreppet kommer att hittas.  
Om Du vill använda platshållare, använder Du SQL-platshållare eller de allmänna platshållarna% eller * för valfritt antal tecken och _ eller? för exakt ett tecken.  
Ett & används automatiskt efter sökbegreppet.  
Använda filter  
En undermeny öppnas med namnen på alla datafält.  
Ett av datafältnamnen är markerat.  
Välj namnet på datafältet där du vill göra sökningen.  
I tabellen visas nu enbart de dataposter som motsvarar sökvillkoret.  
Med ikonen Standardfilter öppnar du dialogen Filter.  
Här kan du filtrera data genom en kombination av flera kriterier  
Med ikonen Ta bort filter sätter du tillbaka vyn till "alla dataposter".  
Radera en datapost  
Klicka på radhuvudet framför den datapost som ska raderas.  
Öppna snabbmenyn och välj kommandot Radera rader.  
Dataposten raderas direkt utan någon fråga.  
Välja kolumntilldelning och datakälla  
På objektlisten finns följande kommandoknappar:  
Kolumntilldelning  
Öppnar dialogrutan Kolumntilldelning för tabell.  
Om du använder en annan datakälla kan du här tilldela datakällans fältnamn fältnamnen som används i %PRODUCTNAME och tvärtom.  
Datakälla  
Öppnar dialogrutan Urval av datakälla där du kan välja datakällan som används för litteraturdatabasen.  
Alla datakällor som är registrerade i %PRODUCTNAME visas.  
Skala  
Med den här funktionen kan du ändra skalan för den visade sidan.  
Med andra procenttal förstorar eller förminskar du vyn.  
Den valda skalan visas på statuslisten.  
Om du använder %PRODUCTNAME -dokument i olika operativsystem märker du kanske att 100% på samma bildskärm och med samma upplösning ser mindre ut med Unix än med Windows.  
Detta beror delvis på att dokument automatiskt förstoras i Windows med cirka 30% för att små teckensnitt ska bli lättare att läsa.  
I Windows måste du alltså ställa in skalan till 75% för att det ska se likadant ut som i andra operativsystem.  
Därför kan ett 8 punkters teckensnitt i en dialogruta se helt annorlunda ut än 8 punkters teckensnitt i ett dokument.  
Zoomfaktor  
Välj någon av de förinställda värdena för förstoring respektive förminskning.  
Hela sidan  
Dokumentsidan visas fullständigt i dokumentfönstret.  
Sidbredd  
Dokumentsidan förstoras respektive förminskas tills även papperskanterna på dokumentet är synliga i fönstret.  
Optimal  
Det här alternativfältet är bara aktivt om Du har markerat ett området.  
Om Du klickar på fältet när Du har markerat ett område förstoras eller förminskas det markerade området så mycket att hela markeringen syns.  
Dokumentsidan förstoras respektive förminskas tills textraden i dokumentet är helt synlig.  
200%  
Med detta alternativ förstoras visningen av dokumentsidan till 200%  
150%  
Här är förstoringen 150%.  
100%  
Här visas sidan i normal storlek.  
75%  
Med detta alternativ förminskas visningen av dokumentsidan till 75% av originalstorleken.  
50%  
Här är förminskningen 50%.  
Steglös  
Här ställer Du in en steglös förstoring eller förminskning.  
Om Du väljer det här alternativet och inte gör någon ändring i rotationsfältet används det senast inställda värdet.  
Du kan också ställa in ett värde i procent med hjälp av pilknapparna bredvid rotationsfältet.  
Funktionslist  
Med det här menykommandot visar eller döljer du funktionslisten.  
Objektlisten  
Det här kommandot visar och döljer Du objektlisten, som innehåller olika sammanhangsberoende funktioner.  
Objektlistens utseende beror på såväl dokumenttyp som den objekttyp som har markerats i dokumentet.  
För vissa typer av arbeten visas flera objektlister samtidigt (t.ex. för tabeller i textdokument).  
Du växlar mellan dem med en liten pilknapp i listens högerkant eller tillhörande snabbmeny.  
När du lämnar ett arbetsområde (t.ex. en tabell) i textdokumentet, registrerar %PRODUCTNAME Writer vilken objektlist som var aktiv, och när du återvänder till det området visas den igen.  
Verktygslist  
Den innehåller olika funktioner som du kan använda i det aktuella dokumentet.  
Verktygslistens innehåll beror på vilken typ av dokument du arbetar med.  
Verktygslisten i ett textdokument skiljer sig t.ex. markant från den i ett tabelldokument.  
Verktygslistens innehåll beror på vilken typ av dokument du arbetar med.  
Verktygslisten i ett textdokument skiljer sig t.ex. markant från den i ett tabelldokument.  
Statuslisten  
Med detta kommando döljer du respektive visar statuslisten i nedre fönsterkanten.  
På statuslisten visas informationen som är definierad under Verktyg - Anpassa - Statuslist.  
Här visas också statusinformation för vissa processer.  
Hela bildskärmen  
Med den här funktionen växlar du mellan helskärm och normalvy.  
Om du vill växla tillbaka till normalvyn kan du använda Kommando Ctrl +Skift+J.  
När du har aktiverat funktionen Hela bildskärmen kan du fortfarande använda de normala tangentkombinationerna för Windows, även om du inte ser menyerna.  
Med kommandot Alt+S kommer du alltså fortfarande till menyn Visa.  
Alla vanliga tangentkombinationer, t.ex. den som du använder när du vill avsluta programmet, går även att använda i helskärmsläge.  
Bekräfta radering  
I den här dialogrutan uppmanas du att bekräfta filåtgärder som kan innebära vissa risker, som när du väljer att Radera filer.  
Du kan antingen bekräfta åtgärden för den aktuella filen eller för alla filer, avvisa åtgärden för den aktuella filen eller avbryta för resterande filer.  
Radera  
Med den här kommandoknappen bekräftar du åtgärden för den aktuella filen.  
Radera alla  
Med den här kommandoknappen bekräftar du åtgärden för den aktuella filen och alla andra markerade filer.  
Radera inte  
Med den här kommandoknappen avvisar Du åtgärden för den aktuella filen.  
Avbryt  
Med den här kommandoknappen avbryter Du åtgärden för den aktuella filen och alla andra filer.  
Färglisten  
På färglisten ser du färgerna på den aktuella färgpaletten.  
Med färglisten kan du välja färg utan att behöva öppna någon dialogruta.  
Klicka på den färg som du vill ge det markerade objektet.  
Om du klickar på färgen som du vill använda med vänster musknapp tilldelas objektet en ny fyllningsfärg.  
Om du klickar med höger musknapp tilldelas objektet en ny linjefärg.  
Du kan också tilldela färgen Osynlig genom att klicka på ikonen uppe till vänster på färglisten.  
Du kan dra färger från färglisten direkt till ritobjekt.  
Om du vill ändra fyllnings - eller linjefärgen låter du färgen falla över ytan eller kanten.  
Om du håller på med att skriva in text i en textram, kan du tilldela en markerad text en ny färg genom att klicka på en färg på färglisten.  
Om du håller på med att skriva in text i en textram, kan du tilldela en markerad text en ny färg genom att klicka på en färg på färglisten.  
Det förankringsbara fönstret på färglisten kan du låta vara öppet medan du redigerar dokumentet.  
Du kan växla mellan färglisten som en förankrad symbollist eller som ett fritt fönster genom att hålla ner Kommando Ctrl -tangenten och dubbelklicka någonstans på ett grått område på listen.  
Om färglisten är ett fönster kan du ändra bredd och höjd.  
Du kan ändra färgerna som visas genom att välja Format - Yta... och klicka på fliken Färger.  
Där kan du ladda en annan färgpalett eller skapa egna färgpaletter som du sparar som filer.  
Symbollister  
Här bestämmer du vilka av symbollisterna som ska visas.  
Med kommandot Redigera kan du förändra symbollisterna.  
Redigera  
Infoga anteckning  
Med den här funktionen infogar du en anteckning vid markörens position.  
Anteckningar är kommentarer som du kan visa och dölja efter egna önskemål.  
Om du redan har infogat och markerat en anteckning heter den här dialogrutan Redigera anteckning.  
Den infogade anteckningen indikeras med en liten gul rektangel i textområdet.  
Dialogrutan Infoga anteckning visas.  
Där kan du läsa och redigera innehållet i anteckningen.  
Utseendet på dialogrutan Redigera anteckning skiljer sig från dialogrutan Infoga anteckning genom två kommandoknappar, med vilka du kan hoppa mellan föregående respektive följande anteckning i dokumentet.  
De knapparna syns bara om du har skapat minst två anteckningar.  
Om du vill kan du inkludera anteckningarna vid utskrift, antingen längst ned på sidan eller sist i dokumentet.  
Den här inställningen gör du under Arkiv - Skriv ut - Fler.  
När du infogar en anteckning i ett tabelldokument ser du inte någon dialogruta utan en förklaringsruta, där du kan skriva texten.  
Klicka utanför rutan när du vill dölja den.  
Infogade anteckningar i tabelldokumentceller indikeras med en röd kvadrat i cellens överkant.  
När du vill läsa texten pekar du med muspekaren på cellen.  
Anteckningen visas som ett hjälptips, och därför måste du ha aktiverat den funktionen på menyn Hjälp - Tips.  
Om du vill redigera anteckningen, klickar du i den cell där den finns och ger sedan återigen kommandot Infoga - Anteckning.  
Om du raderar all text, raderas även anteckningen och dess markeringsruta.  
De visas då på en egen sida efter tabellinnehållet.  
Visa alternativen för tabelldokument genom att välja Format - Sida - Tabell.  
Vid export av dokumentet till en HTML-sida indikeras anteckningarna med <!- - Kommentarer -->.  
Innehåll  
Här kan Du ange information om författaren och skriva en anteckning i textfältet.  
Författare  
Här visas författarens användarinitialer och aktuellt datum.  
Text  
Här skriver Du själva anteckningstexten.  
Skapad av  
Med den här kommandoknappen infogar Du de användarinitialer som anges intill Författare i fältet Text samt aktuellt datum och klockslag.  
Skanna  
Här visas en undermeny med kommandon för skanning av bilder.  
Förutsättningen är du har installerat en skannerdrivrutin.  
För Unix installerar du SANE-paketet, som finns på adressen http: / /www.mostang.com / sane /.  
SANE-paketet måste använda samma libc som %PRODUCTNAME.  
Välj källa  
Rekvirera  
Välj källa  
Med detta kommando öppnar du en dialogruta där du kan välja skanner.  
Välj den skanner som du vill använda.  
Rekvirera  
Med det här kommandot aktiverar du en dialogruta där du styr skanningen.  
Dialogrutan hör till skannerdrivrutinen och är beroende av maskinvaran.  
Mer information om dialogrutan finns i dokumentationen till skannern.  
Specialtecken  
Med den här funktionen kan du infoga ett eller flera specialtecken.  
Du kan öppna den här dialogrutan från de flesta textinmatningsfälten, genom att klicka på Skift + Kommando Ctrl +S.  
Det för tillfället markerade tecknet visas i förstorad form under kommandoknapparna.  
Numret under tecknet motsvarar det numeriska värdet i teckenuppsättningen, som kan vara IBMPC, ANSI, ISO8859-1 eller Mac osv.  
Teckensnitt  
Klicka i kombinationsfältet och välj ett av de installerade teckensnitten.  
När du öppnar dialogrutan från ett textinmatningsfält går det inte att välja något teckensnitt.  
Område  
Välj ett Unicode-område här.  
Tecknen i det valda området visas i teckenurvalsfältet.  
Teckenurvalsfält  
Här ser du de tecken som är tillgängliga i det valda teckensnittet (och i det valda området).  
Välj tecken genom att klicka med musen eller med hjälp av piltangenterna och mellanslagstangenten.  
Tecken  
Här listas i tur och ordning de tecken som du har markerat med musen eller tangentbordet.  
Radera  
Raderar de tecken du markerat utan säkerhetskontroll.  
Hyperlänklisten  
Här kan du sätta på eller stänga av visningen av hyperlänklisten.  
Den är till för redigering och infogning av hyperlänkar och för sökning på Internet.  
Om hyperlänklisten visas, kan du infoga den visade webbadressen på hyperlänklisten i texten med hjälp av ikonen Länk.  
Infoga grafik  
Med den här funktionen infogar du grafik i dokumentet.  
Om du väljer det här kommandot när du har markerat ett grafikobjekt, visas dialogrutan Format - Grafik.  
Under fliken Grafik kan du välja en annan grafikfil som ska ersätta det markerade grafikobjektet.  
Parametrarna (t.ex. Inramning, Hyperlänkar) för det markerade grafikobjektet ändras inte.  
Med det här kommandot (eller ikonen Infoga grafik på verktygslistens utrullningslist Infoga) kommer du till en dialogruta som i stort sett motsvarar dialogrutan Öppna.  
Stil  
Här väljer du en ramformatmall som grafikobjektet infogas med.  
Länka  
Om du markerar den här rutan integreras grafikobjektet inte i dokumentet utan infogas som länk.  
I dokumentet finns då bara en hänvisning till grafikfilen.  
Förhandsvisning  
Du markerar den här rutan om du vill se en förhandsvisning.  
Objekt  
Det här menyalternativet har en undermeny med kommandon som du använder när du vill infoga objekt i ett dokument.  
Du kan välja följande kommandon:  
OLE-objekt  
Ljud  
Video  
Applet  
Formel  
Diagram  
Infoga OLE-objekt  
Med den här funktionen väljer du ut ett OLE-objekt som ska integreras i dokumentet.  
OLE -objekt är objekt som kan länkas med ett måldokument eller integreras.  
De OLE-objekt som hör till dokumentet sparas i minnet så att det ska gå snabbare att ladda dokumentet.  
Det maximala antalet objekt i minnet väljer du under Verktyg - Alternativ - %PRODUCTNAME - Arbetsminne.  
Du kan inte heller dra och släppa dem.  
I andra riktningen kan OLE-objekt integreras i %PRODUCTNAME, men då försvinner länkarna.  
Detta innebär att du kan redigera objekten genom att dubbelklicka på dem men de uppdateras inte när källan ändras.  
Inaktiva OLE-objekt visas transparenta i %PRODUCTNAME Writer.  
Skapa nytt  
På den här sidan definierar du objekttypen för det nya objektet som ska infogas.  
Objekttyp  
Välj objekttypen i den här listrutan.  
Skapa från fil  
Markera det här alternativet om du vill infoga en fil som ett objekt i dokumentet.  
Fil  
I det här området markerar du ett objekt från en fil.  
Fil  
Du kan också ange ett filnamn här.  
Genomsök...  
Om du klickar på den här kommandoknappen visas en dialogruta för filurval där du markerar den fil som ska fogas in.  
Infoga plug-in  
Med den här funktionen infogar du en plug-in.  
Fil / URL  
Du kan också ange ett filnamn här.  
Genomsök...  
Om du klickar på den här kommandoknappen visas en dialogruta för filurval där du markerar den fil som ska fogas in.  
Alternativ  
I det här fältet anger du parametrar som ska övertas vid export till ett HTML-dokument.  
Den här funktionen kan du bara använda när du känner till de exakta parametrarna för insticksprogrammet.  
Infoga applet  
Med den här funktionen infogar du ett applet -program.  
Fil  
I det här området finns fält för definition av Klass och Class Location.  
Klass  
I fältet Klass visas applet-klassen, t.ex. "Ticker".  
Class Location  
I det här fältet står klassplaceringen för Applet-programmet, d.v.s. den plats där Applet-programmet är arkiverat.  
Genomsök...  
Genom att klicka på kommandoknappen kan du antingen söka efter klass eller Class Location för Applet-programmet, beroende på i vilket av fälten markören står.  
Alternativ  
I det här fältet anger du parametrar för Applet-programmet.  
Infoga ljud  
Med hjälp av den här funktionen kan du infoga ljud.  
Dialogrutan Infoga ljud motsvarar den dialogruta som du kan öppna med Arkiv - Öppna.  
Välj ut katalogen och namnet på ljudfilen och infoga önskat ljud i dokumentet med kommandoknappen Infoga.  
Infoga video  
Med den här funktionen infogar du en video.  
Dialogrutan Infoga video motsvarar den dialogruta som du kan öppna med Arkiv - Öppna.  
Välj ut katalogen och namnet på videofilen, och infoga önskad fil i ditt dokument med kommandoknappen Infoga.  
Autoformat diagram  
Här infogar du ett diagram i dokumentet.  
När du klickar på ikonen Infoga diagram ändras markören till ett litet kors med en diagrambild.  
Rektangelns storlek visar hur stort diagrammet blir.  
Du kan även ändra diagrammets storlek och läge senare.  
Då tillåts också multipel markering.  
Mer information om multipel markering med luckor finns i exemplet.  
Det markerade området anges i textfältet Område i dialogrutan Autoformat Diagram (1-4).  
Klicka på ikonen till höger om fältet Område.  
I förhandsvisningen i dialogrutan Autoformat Diagram visas de data som du har markerat i tabellen.  
Antalet datapunkter som visas är begränsat till 20 för att visningen inte ska ta för lång tid.  
Av samma skäl är det inte säkert att du genast ser designändringar i ett diagram i förhandsvisningen.  
Om det redan finns ett diagram i tabelldokumentet och du vill ändra dataområdet markerar du bara det nya området och drar det till diagrammet med musen.  
Då visas dialogrutan Ändra källdataområde där du kan definiera etiketten för det nya diagrammet.  
Du kan också ändra dataområdet via snabbmenyn.  
Med kommandot Ändra dataområdet... visar Du dialogrutan Ändra diagramdataområdet.  
Denna är uppbyggd på samma sätt som dialogrutan AutoFormat Diagram - Sidan 1 av 4.  
Här ändrar Du dataområdet.  
Med menykommandot Infoga - Objekt - Diagram eller ikonen Infoga diagram som finns på utrullningslisten Infoga objekt öppnar du dialogrutan Autoformat Diagram (1-4).  
Sidorna 2 till 4 är identiska med sidorna 1 till 3 i motsvarande dialog som visas när du har markerat ett diagram och väljer kommandot Format - AutoFormat.  
Autoformat Diagram - Sidan 1 av 4  
Urval  
I detta område väljer Du ut vilka celler i tabellen som ska användas i diagrammet.  
Område  
Definiera här det tabellområde som Du vill skapa ett diagram för.  
Cellen under B1 heter B2 osv.  
Så här anger Du ett tabellområde:  
Ange först den cell som är överst till vänster.  
Skriv in ett kolon (:) och ange cellen längst ned till höger.  
Om Du vill ange ett område som sträcker sig från den första cellen överst till vänster till cellen i tredje raden och tredje kolumnen skriver Du så här:  
A1:C3.  
Då övertas området automatiskt.  
I tabelldokument markeras ett sammanhängande område med värden automatiskt när du klickar på ikonen Diagram, under förutsättning att du har placerat cellmarkören i området.  
Första raden som etikett  
Markera den här rutan om du har markerat kolumnöverskrifterna i den första raden i området.  
De används då som etiketter i diagrammet.  
Första kolumnen som etikett  
Markera den här rutan om du har markerat radöverskrifterna i den första kolumnen i området.  
De används då som etiketter i diagrammet.  
Utdata i tabell  
Om Du vill infoga ett diagram i ett %PRODUCTNAME Calc-dokument som består av flera tabeller anger Du i denna listruta i vilken tabell diagrammet ska infogas.  
<< Tillbaka  
I dialogrutan kan Du visa de val som Du har gjort på föregående sida.  
Aktuella inställningar bibehålls.  
Denna knapp är endast tillgänglig fr o m det andra redigeringssteget.  
Nästa >>  
När Du klickar på den här knappen använder AutoPiloten de aktuella inställningarna i dialogrutan och går vidare till nästa sida.  
Om Du har kommit till den sista sidan i dialogrutan kan knappen inte väljas.  
Färdigställ  
När Du klickar på knappen skapar AutoPiloten ett diagram som infogas i dokumentet utifrån de inställningar som Du har gjort  
Exempel på multimarkering  
Om du markerar ett sammanhängande område av celler och infogar ett diagram används det markerade området för diagramdata.  
Ett försök görs att filtrera bort de rader och kolumner som finns mellan de markerade cellerna och därefter sammanfoga de resterande områdena.  
Om detta går utan luckor skapas diagrammet med de sammanfogade områdena.  
Om det fortfarande finns luckor kvar kommer de enskilda markeringarna att skrivas under varandra.  
Anta att du har gjort följande markering:  
Här skapas automatiskt ett diagram för januari, februari, mars, april och maj för Hylla 1.  
Titta på följande multimarkering:  
Diagrammet kommer inte att säga så mycket.  
Nu tar vi en multimarkering som kan sammanfogas:  
Här skapas ett diagram för februari och mars, för hylla 2 och 4.  
Men varför ska du markera den tomma cellen A1?  
Försök utan A1:  
Den här multimarkeringen fungerar också!  
Du skapar ett diagram för februari och april, för hylla 2 och 4.  
Autoformat Diagram - sida 1 av 3 Autoformat Diagram - sida 2 av 4  
På den här sidan i dialogrutan Autoformat Diagram väljer du diagramtyp.  
Förhandsvisning  
Här kan du se hur den diagramtyp som du har skapat kommer att se ut.  
Förhandsvisningen förekommer även på de andra sidorna.  
Visa textobjekt i förhandsvisning  
Markera den här rutan om du vill visa textobjekt, t.ex. förklaringar, överskrifter och axelrubriker, med diagramtypen i förhandsvisningsfältet.  
Fältet syns också på de andra sidorna.  
Dataserier i:  
Rader  
Kolumner  
Välj en diagramtyp  
Här väljer Du önskad diagramtyp.  
Fortsätt till Autoformat Diagram - sida 2 av 3 Mera om Autoformat Diagram - sida 3 av 4  
Autoformat Diagram - sida 2 av 3 Autoformat Diagram - sida 3 av 4  
Här kan du bestämma hur dina diagram ska visas.  
Dataserier i:  
Rader  
Kolumner  
Välj ut en variant  
Här kan du välja den variant du föredrar.  
Mer information om varianterna finns här.  
Gitterlinjer  
I det här området kan Du lägga in gitterlinjer som bakgrund i den diagramtyp som Du har valt.  
X-axel  
Om Du vill att gitterlinjerna ska utgå från x-axeln klickar Du här.  
Y-axel  
Om Du vill att gitterlinjerna ska utgå från y-axeln klickar Du här.  
Z-axel  
Om Du vill att gitterlinjerna ska utgå från z-axeln klickar Du här.  
Detta alternativ finns förstås bara för tredimensionella diagram.  
Fortsättning på Autoformat Diagram - sida 3 av 3 FortsÃ¤ttning pÃ¥ Autoformat Diagram - sida 4 av 4  
AutoFormat Diagram - sidan 3 av 3 AutoFormat Diagram - sidan 4 av 4  
På den här sidan definierar du bland annat en rubrik för diagrammet.  
Diagramrubrik  
Här definierar du om diagrammet ska tilldelas ett namn.  
I textfältet anger du en diagramrubrik.  
Dataserier i  
I detta område väljer du om dataserierna ska visas i rader eller kolumner.  
Rader  
Markera det här alternativfältet om du vill att dataserierna ska visas i rader.  
Kolumner  
Markera det här alternativfältet om du vill att dataserierna ska visas i kolumner.  
Detta är standardinställningen i %PRODUCTNAME.  
Förklaring  
Klicka här om diagrammet ska ha en förklaring.  
Axelrubrik  
I det här området tilldelar du varje axel en rubrik.  
X-axel  
Här tilldelar du X-axeln (den vågräta axeln) en rubrik.  
Y-axel  
Här ger du Y-axeln (den lodräta axeln) en rubrik.  
Z-axel  
Här anger du en rubrik för Z-axeln.  
Det går bara att välja det här alternativet för tredimensionella diagram.  
Ändra källdataområde  
Etikett  
Här anger du om du vill använda den första kolumnen och första raden i det markerade området som etikett för diagrammet.  
Markera den här rutan om du har markerat radöverskrifterna i områdets första kolumn.  
De övertas då som etikett i diagrammet.  
Markera den här rutan om du har markerat kolumnöverskrifterna på områdets första rad.  
De övertas som etikett i diagrammet.  
Formel  
Med den här funktionen startar du formel-editorn %PRODUCTNAME Math som anvÃ¤nds till att infoga matematiska formler.  
När du väljer det här kommandot visas fönstren Kommandon och Urval där du kan välja formel -kommandon.  
Men du kan även skriva en text direkt i textdokumentet, markera texten och sedan välja menyn Infoga - Objekt - Formel.  
Det markerade innehållet används som formel.  
Infoga ram  
Med den här funktionen infogar du en ram i dokumentet.  
Om du vill skapa HTML-sidor med flytande ramar, ställer du in exportalternativet "MS Internet Explorer 4.0" under Verktyg - Alternativ - Ladda / spara - HTML-kompabilitet.  
Den flytande ramen förses med taggarna <IFRAME> och < / IFRAME>.  
De här taggarna kan inte utvärderas av alla webbläsare.  
Definiera egenskaperna för ramen som du vill infoga i dialogrutan Ram - egenskaper.  
Datakällor  
Här sätter du på och stänger av datakällvyn.  
Databaslisten med särskilda styrelement för datavisningen visas.  
Kommandot Datakällor på menyn Visa är bara tillgängligt när ett text - eller tabelldokument är öppet.  
För text - och tabelldokument med formulärfunktioner via Kontrollfält med databaskoppling.  
På objektlisten för datavyn visas ikoner för sortering och filtrering av datavisningen samt andra sammanhangsberoende ikoner.  
Kommandoelementen i datavyns undre kant används för att navigera i de visade dataposterna.  
Grafik  
Här väljer du från vilken källa du vill infoga grafik.  
Från fil  
Standard  
Med det här kommandot återställer du ändringar i den markerade dataseriens datapunkter till deras ursprungliga formatering.  
Med det här kommandot formaterar du om det markerade stycket med motsvarande styckeformat.  
Med det här kommandot återställer du de markerade cellerna till standardformatet.  
Med det här kommandot formaterar du om det markerade objektet med motsvarande format.  
Den nya formateringen orienterar sig efter formatmallarna.  
När du skriver en ny text i ett stycke och har försett texten med direkta format men vill fortsätta att skriva utan direkt formatering trycker du bara en gång på höger piltangent.  
Då skriver du vidare med samma format som det första tecknet i stycket har.  
Använd Format - Standard om du vill omvandla en hyperlänk i en text i en tabell till normal text igen.  
Markera då cellområdet med länken och formatera den med standardformatet.  
Markera länken, eventuellt med tecknen före och efter, eller med Alternativ Alt -tangenten nedtryckt.  
Kommandot finns också på snabbmenyn.  
Tecken  
Med den här funktionen kan du bland annat ställa in teckensnitt och teckeneffekt.  
Dessutom kan du tilldela tecknen en hyperlänk eller ett makro.  
Teckensnitt  
Hyperlänk  
Tecken Teckensnitt  
Här finns funktioner för redigering av teckensnitt, teckenstil, teckenstorlek, språk och teckenfärg.  
Om markören står inuti ett ord, används funktionen på hela ordet.  
Om ett område är markerat, gäller den hela området.  
Om inget området är markerat, används den nya funktionen vid skrivning av text från markörens plats.  
Du ser följande områden:  
Teckensnitt för västlig text - välj inställningarna för västlig text här, t.ex. i latinska teckenuppsättningar.  
Teckensnitt för asiatisk text - välj inställningarna för asiatisk text här, t.ex. i kinesiska, japanska och koreanska teckenuppsättningar.  
Teckensnitt  
Här kan du skriva eller välja namnet på ett teckensnitt.  
Teckenstil  
Här kan du ange eller välja en stil.  
Även för detta finns ikoner på objektlisten.  
Teckenstorlek  
Här kan du ange eller välja ut en teckenstorlek.  
För fritt skalbara teckensnitt kan du även ange mellanstorlekar.  
När du redigerar mallar som baserar på överordnade mallar kan du ändra teckenstorleken.  
Du kan ange storleken i procent (t.ex. 150% eller 50%) eller som skillnad mätt i punkter (t.ex. -2pt eller +5pt).  
Språk  
Här bestämmer du vilket språk som ska användas vid rättstavningskontrollen.  
Den här möjligheten finns bara i dialogrutan Format - Cell - Tal, däremot inte (för textobjekt) i dialogrutan Format - Tecken - Teckensnitt.  
Språkmodulerna som är installerade i ditt %PRODUCTNAME är markerade med en bock.  
Teckenfärg  
Här väljer du teckenfärg.  
Om rutan Svart utskrift är markerad i dialogrutan Verktyg - Alternativ - Textdokument - Skriv ut, kommer färgändringar i texten inte att skrivas ut.  
Välj Automatiskt om färgen som är inställd i systemet ska väljas som teckenfärg.  
Om du vill definiera egna färger, stänger du dialogrutan och väljer i dialogrutan Verktyg - Alternativ - %PRODUCTNAME - Färger en färgvariation i färgtabellen.  
Redigera den, ge den ett nytt namn och klicka på Lägg till.  
Nu kan du välja den nya färgen sist i kombinationsfältet Färg.  
Om du klickar länge på ikonen öppnas en utrullningslist där du kan välja en textfärg.  
Om du klickar kort på ikonen tilldelar du den markerade texten färgen som du har valt eller så aktiveras symbolen för färgöverstrykning.  
Om symbolen för färgöverstrykning (färgburken) eller tilldelningsläge är aktiverad kan du ångra genom att klicka en gång med den högra musknappen någonstans i dokumentet.  
Den här funktionen har du nytta av om du vill upphäva den senaste tilldelningen med symbolen för färgöverstrykning (färgburken) eller tilldelningsläge.  
Men du kan också ångra andra steg av misstag om du inte ser upp med var du klickar.  
Om ett felmeddelande visas när du startar %PRODUCTNAME med information om att vissa teckenuppsättningar i %PRODUCTNAME inte kan hittas, kan du i efterhand skapa dem med hjälp av setupprogrammet i reparationsläge.  
Teckeneffekt  
Här kan du välja teckeneffekter.  
Understrykning  
Välj typ av understrykning.  
Även mellanrum och tabbar stryks under om du markerar rutan Ordvis.  
När bara upphöjd text stryks under blir även understrykningen upphöjd.  
När upphöjd text stryks under tillsammans med normal text stannar understrykningen kvar på baslinjen.  
Färg  
Här väljer du färg för understrykningen.  
Effekter  
I det här området kan du välja en effekt i kombinationsfältet och markera rutorna Kontur, Skugga och Blinkande en och en eller tillsammans.  
Effekter  
Välj mellan följande effekter:  
(Utan) - återställer en tilldelning av en effekt.  
Versaler - tecknen visas med stora bokstäver (inte omvandlade).  
Gemener - tecknen visas med små bokstäver (inte omvandlade).  
Titel - den första bokstaven i varje ord visas som stor bokstav.  
Kapitäler - alla tecken visas med stora bokstäver.  
Vid ord som börjar med en stor bokstav är den första bokstaven något större än bokstäverna som kommer efter.  
Genomstrykning  
Välj typ av genomstrykning.  
Vid export till MS Word-format ignoreras alla genomstrykningar utom enkel genomstrykning, d.v.s. de visas som enkla genomstrykningar eftersom Word inte klarar andra typer.  
Ordvis  
Om den här rutan är markerad avbryts under - eller genomstrykning avbryts i mellanrummen mellan orden.  
Kontur  
Om du markerar här visas bara tecknens konturer.  
Den här effekten går inte använda på alla teckensnitt.  
Skugga  
Här har du möjlighet att förse tecknen med skugga.  
Blinkande  
När du markerar den här kryssrutan visas markerad text som blinkande.  
Det går inte att ställa in blinkfrekvensen.  
Betoningstecken  
Välj betoningstecken här.  
Position  
Över text eller Under text.  
Relief  
Välj här bland effekterna (Utan), Upphöjt eller Graverat.  
Tal / format  
Här definierar du formaten för visning av tal.  
Kategori  
Här visas de olika kategorierna för alla format.  
Speciella egenskaper för talformat  
När du räknar med valutor i en tabell används valutaformatet från den formaterade cellen.  
Detta gäller också för de grundläggande räkneoperationerna.  
Du kan tilldela cellerna ett annat format manuellt.  
Format  
Här finns en förteckning över alla definierade format för en bestämd kategori.  
Det som Du markerar i denna listruta avgör vilka poster som visas i fältet Formatbeskrivning och om området Alternativ är aktiverat.  
Listrutan Kategori Valuta  
Speciella egenskaper för talformat  
I detta visningsfält finns många valutor att välja mellan (t ex Euro).  
För varje valuta finns dessutom flera format.  
Valutasymbolen visas också.  
Valutaformatet kan du ställa in oberoende av språk eller land.  
Formatkoden är uppbyggd enligt formatet [$xxx-nnn].  
För Sverige och kronan ställs alltså [$kr-41D] in.  
Talet är en programintern landsidentifierare som du inte behöver ange om du vill definiera egna format.  
Särskilda banksymboler som t.ex. SEK eller EUR kodas alltid utan landsidentifikation.  
När flera valutaformat är definierade för ett språk i ditt operativsystem är valutaformaten som visas i listrutan en kombination av inställningarna i fältet Språk och fältet Format.  
Använd tusentalsavgränsare för att på ett smidigt sätt formatera valutaformat enligt mönstret 00 tkr.  
Om du exempelvis vill skapa alla belopp enligt formatet "tusen kr med en decimal" anger du 0,0 [$tkr] som formatkod.  
1,124 tkr.  
Språk  
I det här kombinationsfältet kan du välja ett annat språk än det förinställda om du vill använda ett utländskt talformat.  
Språkurvalet påverkar datum - och valutaformatet.  
Om du byter språk kommer alla celler som formaterats med standarddatumformat eller med standardvalutaformat att anta det nya landsspecifika datum - eller valutaformatet.  
Detta gäller inte format som du själv har definierat.  
Anta att du har angett "1 kr" i en cell och därefter sparar dokumentet.  
Den här filen öppnas sedan exempelvis i ett engelskt system.  
Standardvalutaformatet kommer inte att användas för cellen och din inmatning bibehålls i systemet på annat språk.  
Källformat  
Om den här rutan är markerad, väljer %PRODUCTNAME talformat från cellformatet för cellerna som diagrammet skapades av.  
Om du vill ha ett eget talformat måste du upphäva markeringen av det här fältet först.  
Alternativ  
Här kan du komplettera visningen av cellinnehållet i egna format.  
Antal decimaler  
Här definierar Du antalet decimaler för tal som ska formateras enligt ett bestämt talformat.  
Inledande nollor  
Här definierar Du antalet inledande nollor.  
Negativa värden i rött  
Markera den här rutan om du vill att negativa tal som formateras i ett visst talformat ska visas i rött.  
Tusentalsavgränsare  
Markera den här rutan om stora tal som formateras enligt ett bestämt talformat ska avgränsas med ett blanksteg.  
Formatbeskrivning  
Här visas formatbeskrivningen som motsvarar det format som Du markerat i listrutan Format.  
Du kan också definiera egna formatbeskrivningar genom att välja "Användardefinierad" i listrutan Kategori.  
För användardefinierade format får Du tillgång till ikonerna Lägg till, Ta bort och Ändra kommentar.  
Lägg till  
Med denna ikon lägger Du till formatbeskrivningen till den användardefinierade kategorin.  
Ta bort  
Med denna ikon tar Du bort formatbeskrivningen för den användardefinierade kategorin.  
Ändringen träder i kraft när Du startar om programmet.  
Ändra kommentar  
Med denna ikon infogar eller ändrar du en kommentar som visas under fältet Formatbeskrivning.  
Som standard står här "Användardefinierad".  
Om du har definierat en egen formatbeskrivning klickar du på den här ikonen.  
En textruta öppnas där du kan skriva en kommentar till det egna formatet.  
Kommentarrad  
Här anger Du en kommentar för Dina egna format.  
När Du klickar på ikonen Ändra kommentar ändras kommentaren.  
Formatkod; talTalformatkoder  
Talformatkoderna (under Format - Cell - Talformat) kan bestå av upp till tre avsnitt som du gränsar av med hjälp av semikolon (;).  
Om en kod innehåller två avsnitt så gäller det första avsnittet för positiva värden och noll och det andra avsnittet för negativa värden.  
Om en kod innehåller tre avsnitt så gäller det första avsnittet för positiva värden, det andra avsnittet för negativa värden och det tredje för noll.  
Du låter då det första avsnittet gälla om det uppfyller det första villkoret, det andra avsnittet om det uppfyller det andra villkoret och det tredje avsnittet utförs om inget av villkoren uppfylls.  
Ett exempel finns längst ned på denna sida.  
Använd Vetenskap för att visa tal vars sifferantal överstiger cellbredden.  
Om Du vill visa ett bestämt antal siffror (0 eller #) till höger och vänster om decimaltecknet infogar Du ett decimaltecken (i Sverige ett kommatecken) i talformatet.  
Om formatet redan innehåller nummertecknet (#) till vänster om decimaltecknet kommer tal som är mindre än 1 att börja med decimaltecknet.  
Använd följande formatkoder i ett avsnitt om Du vill skapa platshållare för tal.  
Om ett tal har fler siffror till höger om decimaltecknet än det finns platshållare för i formatet, avrundas talet till den decimal som motsvarar platshållaren.  
Om talet har fler siffror till vänster om decimaltecknet än det finns platshållare för i formatet, visas dessa.  
Platshållare  
Betydelse  
#  
inga ytterligare nollor visas.  
0 (noll)  
fler nollor visas om talet har färre siffror än det finns nollor i formatet.  
Talformat  
Formatkod  
3456,78 som 3456,8  
####,#  
9,9 som 9,900  
#,000  
13 som 13,0 och 1234,567 som 1234,57  
#,0#  
5,75 som 5 3 / 4 och 6,3 som 6 3 / 10  
#??? /???  
,5 som 0,5  
0,##  
Antalet frågetecken anger hur många siffror täljare och nämnare kan bestå av.  
Bråk som inte passar in, visas som flyttal.  
Infoga en punkt i talformatet om Du vill visa en punkt som tusentalsavgränsare eller om Du vill att ett tal ska visas som en multipel av tusen.  
Talformat  
Formatkod  
15000 som 15.000  
#.###  
16000 som 16  
#.  
Du ställer in färgen för ett avsnitt genom att infoga färgens namn inom hakparenteser.  
CYAN  
GRÖN  
SVART  
BLÅ  
MAGENTA  
RÖD  
VIT  
GUL  
Talformatkoder för datumformat  
Infoga följande formatkoder om du vill visa dagar, månader och år.  
Format  
Formatkod  
Månad som 3.  
M  
Månad som 03.  
MM  
Månad som jan-dec  
MMM  
Månad som januari-december  
MMMM  
Första bokstaven i månadsnamnet  
MMMMM  
Dag som 28.2.  
D  
Dag som 02  
DD  
Dag som må-sö  
NN eller DDD  
Dag som söndag till lördag  
NNN eller DDDD  
Dag med följande skiljetecken, t.ex. som måndag-söndag  
TTTT  
År som 00-99  
JJ  
År som 1900-2078  
JJJJ  
Kalendervecka  
WW  
Kvartal som Q1 till Q4  
Q  
Kvartal som kvartal 1 till kvartal 4  
QQ  
Era i japansk Gengou-kalender, ett tecken långt (möjliga värden:  
M, T, S, H)  
G  
Era, förkortad form  
GG  
Era, fullständigt namn  
GGG  
Årtal i en era, utan inledande nolla vid år som bara består av en siffra  
E  
Årtal i en era, med inledande nolla vid år som bara består av en siffra  
EE eller R  
Era, fullständigt namn och år  
RR eller GGGEE  
Du kan lägga till följande teckensträngar i formatkoderna om du vill använda en viss kalender.  
Om det saknas en fast inmatad kod väljer %PRODUCTNAME bästa möjliga kalender som ska användas.  
[~gregorian]  
Gregoriansk kalender  
[~gengou]  
Japansk Gengou-kalender  
[~ROC]  
Koreansk kalender  
Alla kalenderformat är beroende av "Locale", språkvarianten som du kan välja under Verktyg - Alternativ - Språkinställningar - Språk.  
Ett exempel: datumformatskoden E, EE, R eller RR ställer om kalendern till den första icke-gregorianska kalendern som är registrerad för den aktuella språkvarianten.  
Om du använder en japansk språkvariant är det Gengou-kalendern.  
Om du använder en koreansk språkvariant är det ROC-kalendern.  
Om ingen ytterligare kalender är angiven för språkvarianten används den gregorianska kalendern.  
Om du räknar med cellreferenser där minst en referens har tilldelats ett datum - eller tidsformat visas resultatet automatiskt med lämpligt format.  
Du kan tilldela formelcellen ett annat format manuellt.  
Det finns följande alternativ:  
Utgångsformat  
Resultatformat  
Datum + Datum  
Tal (Dagar)  
Datum + Tal  
Datum  
Datum + Tid  
Datum&Tid  
Datum + Datum&Tid  
Tal  
Tid + Tid  
Tid  
Tid + Tal  
Tid  
Tid + Datum&Tid  
Datum&Tid  
Datum&Tid + Datum&Tid  
Tid  
Datum&Tid + Tal  
Datum&Tid  
Tal + Tal  
Tal  
Datum&Tid-formatet visar både datum och klockslag och skapas så snart Du lägger ihop ett värde i datumformat med ett i tidformat.  
Förutom att addera kan Du förstås subtrahera, multiplicera och dividera värden.  
Standardvärdet är 1899-12-30.  
Anger Du ett årtal med två siffror bestäms med hjälp av 29 / 30-regeln om det betyder 19xx eller 20xx.  
Ett datum som 1.1.30 betyder däremot 1.1.1930.  
När Du öppnar ett %PRODUCTNAME Calc-dokument innan version 5.0 gäller den gamla regeln som säger att (nästan) alla tvåsiffriga årtal får prefixet 19 (förutom eventuellt de senaste dagarna år 1899, se ovan).  
Talformatkoder för tidsformat  
Infoga följande formatkoder om du vill visa timmar, minuter och sekunder.  
Format  
Formatkod  
Timmar som 0-23  
h  
Timmar som 00-23  
hh  
Minuter som 0-59  
m  
Minuter som 00-59  
mm  
Sekunder som 0-59  
s  
Sekunder som 00-59  
ss  
Du kan använda decimaltecknet i formatkoden för att visa delar av sekunder.  
Du kan t.ex. visa tiden 01:02:03,45 med koden hh:mm:ss,oo.  
Om du vill visa tid som är längre än 24 timmar eller mer än 60 minuter eller sekunder sätter du den yttersta vänstra delen av tidskoden inom hakparentes.  
Exempelvis visar tidskoden [h ]:mm:ss mer än 24 timmar.  
Du kan också räkna med tidsformaten.  
Detta är t.ex. praktiskt vid subtraktioner enligt mönstret: tid=sluttid-starttid.  
Om Du skriver in ett klockslag som 02:03,45, 01:02:03,45 eller 25:01:02 tilldelas följande format såvida Du inte redan har angett ett annat tidsformat:  
MM:SS,00, [HH]:MM:SS,00 eller [HH ]:MM:SS.  
Vid addition och subtraktion av tider visas värdet i en formelcell i ett motsvarande format, beroende på resultatet.  
Detta är t ex praktiskt vid beräkning enligt mönstret = sluttid-starttid eller =( sluttid-starttid )*24*timlön.  
Talformatkoder för valutaformat  
Det valutatecken som är tillgängligt enligt språkvarianten är förvalt som standard för valutaformatet om du har valt standard som språk.  
Eurovalutan infogar du med en av följande formatkoder:  
#.##0,00 "EUR" ;[RED]-#.##0,00 "EUR"  
#.##0,00 [$€-407] ;[RED]-#.##0,00 [$€-407]  
Banksymbolen EUR är den internationella förkortningen för euro.  
Det andra exemplet visas om du väljer posten "€tyska (Tyskland)" i kombinationsfältet Format.  
Delen [$€-407] av formatkoden betyder att eurotecknet (€) och språkvarianten 407 används.  
Du väljer koden för en språkvariant i kombinationsfältet Format.  
Koden registreras då automatiskt korrekt i fältet Formatbeskrivning.  
Talformatkoder för text och blanksteg  
Om Du vill visa tecken sätter Du dem antingen inom dubbla citattecken eller placerar ett omvänt snedstreck (\) framför dem.  
Om Du vill skapa ett blanksteg med samma bredd som ett tecken i ett talformat infogar Du ett understreck (_) följt av tecknet.  
Om du skriver ett understreck och en slutparentes visas exempelvis positiva tal och negativa tal justerade till varandra i parenteser.  
Om Du vill innefatta ett textavsnitt i ett talformat infogar Du @-tecknet i talformatet.  
Text som Du har angett i en cell formateras enligt det avsnitt som innehåller @-tecknet.  
Om det inte finns något textavsnitt i formatet påverkas inte den text som Du skriver av formatet.  
Ytterligare talformatkoder  
Då multipliceras talet med 100 och procenttecknet läggs till.  
Vetenskapsformat  
Om Du vill visa tal i formatet Vetenskap infogar Du följande formatkod i ett avsnitt.  
Om formatet innehåller 0 eller #-tecknet till höger om E-, E+, e - eller e + visas talet i ett tabelldokument i formatet Vetenskap och "E" eller "e "infogas.  
Antalet nollor eller #-tecken till höger bestämmer antalet siffror i exponenten.  
Med E - eller e - visas ett minustecken vid negativa exponenter.  
Med E + eller e + visas ett minustecken vid negativa exponenter och ett plustecken vid positiva exponenter.  
Format med prefix och suffix  
Du kan utöka talformaten med text före och efter (prefix och suffix) och formatera celler med denna kod.  
Definiera t.ex. följande formatkod:  
0 "plus";0 "minus";0 "noll"  
Dessutom följs de som suffix av texten inom citattecken (texten visas utan citattecken i cellerna).  
Om Du t ex anger "1" i en cell blir resultatet "1 plus ".  
Om Du anger "-5" får Du resultatet "5 minus ".  
Villkor i talformaten  
Du kan lägga in villkor för jämförelse med tal direkt i formatkoden.  
Här följer ett exempel.  
###[ <=4][GRÖN]#.##0,00 ;[>7][RÖD]#.##0,00 ;[BLÅ ]#.##0,00  
Här formateras en cell enligt talformatet #.##0,00.  
Vid ett värde över 7 blir den röd.  
I övriga fall är textfärgen blå.  
Du kan använda relationsoperatorerna <, <=, >, >=, = och <> tillsammans med valfria tal.  
Landsspecifika talformat  
I dialogrutan Talformat Under fliken Tal kan du använda landsspecifika formatdefinitioner.  
Både standard-datumformatet och standard-valutaformatet administreras landsspecifikt av %PRODUCTNAME.  
Valutaformaten i %PRODUCTNAME kan ställas in oberoende av land resp. språk.  
Du kan också definiera egna valutaformat i %PRODUCTNAME.  
Men när du använder dem måste du tänka på att export av data inte sker oberoende av operativsystem.  
Dessutom har du tillgång till valutaformatet euro i %PRODUCTNAME.  
Hyperlänk  
Här kan du tilldela de markerade tecknen en hyperlänk.  
En hyperlänk, ofta kallad "länk", är en hänvisning till ett dokument på Internet eller i det lokala systemet.  
Du kan också ange ett HTML-ankare som har infogats som bokmärke, om du vill hänvisa till en viss plats i det angivna dokumentet.  
En annan möjlighet att ange och redigera hyperlänkar finns i hyperlänkdialogen.  
Hyperlänk  
I det här området väljer du måldokument och målram.  
URL  
I det här fältet anger Du måldokumentets fullständiga webbadress, som ska laddas när man klickar på hyperlänken.  
Måldokumentet ersätter det aktuella dokumentet, om Du inte anger en annan målram (Ram).  
Om du vill ändra en URL som redan står i texten kan du bara skriva över den i dokumentet.  
Välj ut...  
Via den här kommandoknappen kommer Du till dialogrutan Öppna.  
Välj en målfil i filsystemet eller på en FTP-server på Internet.  
Tips!  
Här skriver Du den text som ska visas som namn på hyperlänken i dokumentet.  
Händelser...  
Med den här kommandoknappen öppnar du dialogrutan Tilldela makro.  
Här kan du tilldela hyperlänken ett makro som ska utföras.  
Namn  
I det här textfältet kan du tilldela hyperlänken ett ankarnamn.  
En NAME-tagg infogas på följande sätt:  
<A HREF=" http: / /www.sun.com / "NAME="Namntext" TARGET="_blank ">Hänvisningstext< / A>  
Du kan nu hoppa till den här hyperlänken från en annan plats.  
NAME-taggen fungerar bara i HTML-dokument.  
Ram  
I det här kombinationsfältet väljer du bland de givna alternativen den målram där måldokumentet ska visas.  
Om du inte anger någon målram, ersätts det aktuella dokumentet av måldokumentet.  
Teckenformatmallar  
I det här området väljer du teckenformatmallar till den aktuella hyperlänken.  
En använd länk markeras på annat sätt.  
Använd länk  
Här väljer du teckenformatmall till den aktuella hyperlänken om den redan har använts.  
Oanvänd länk  
Här väljer du teckenformatmall till den aktuella länken om den ännu inte har använts.  
Teckenposition Position  
Här bestämmer du position och avstånd för tecknen.  
Position  
Här bestämmer du position för tecknen uppåt eller neråt.  
Upphöjd  
Du kan välja en förminskning.  
Normal  
Tecknen återges i den aktuella teckenstorleken på textbaslinjen.  
Nedsänkt  
Med det här alternativet återges tecknen med en nedsänkt position.  
Du kan välja en förminskning.  
Höj / sänk med  
Här definierar du den relativa placeringen av den upphöjda eller nedsänkta texten i relation till den aktuella teckenstorleken.  
Rel. teckenstorlek  
Här definierar du den relativa storleken på den upphöjda eller nedsänkta texten i relation till den aktuella teckenstorleken.  
Automatiskt  
Om du väljer den här funktionen görs den relativa placeringen av den upphöjda eller nedsänkta texten automatiskt.  
Avstånd  
Här ändrar du avståndet mellan de enskilda tecknen.  
Avstånd  
Här definierar du avståndet mellan tecknen.  
Standard - väljer det teckenavstånd som har definierats i teckensnittet  
Spärrat - en förstoring av teckenavståndet  
Smalt - en förminskning av teckenavståndet  
Avståndet infogas före tecknen.  
Du kan ändra avståndet mellan två bokstäver genom att tilldela den första bokstaven en spärrad eller smal stil.  
Avstånd med  
Här definierar du avståndet i den typografiska måttenheten punkt.  
Parvis kerning  
Markera den här rutan om teckenavståndet ska anpassas automatiskt för vissa bokstavskombinationer.  
För att det ska gå att använda parvis kerning i %PRODUCTNAME måste din skrivare och skrivardrivrutin ha stöd för det.  
Dessutom måste kerningpar vara definierade i det använda teckensnittet.  
Rotation / skalning  
Här väljer du rotationsvinkeln för tecken.  
0 grad  
Det här alternativet bestämmer justeringen från vänster till höger.  
90 grader  
Med det här alternativet roterar du tecknen 90 grader moturs.  
270 grader  
Med det här alternativet roterar du tecknen 270 grader moturs.  
Anpassa till rad  
Välj här så anpassas tecknen till raden.  
Skala bredd  
Välj här den procentuella skalningen av bredden.  
Asiatisk layout  
Här definierar du inställningarna för dubbla rader i asiatisk layout.  
Markera först tecknen som du vill skriva på dubbla rader i dokumentet och använd sedan den här funktionen.  
Dubbla rader  
Här väljer du om du vill skriva de markerade tecknen på dubbla rader.  
Skriva på dubbla rader  
Markera den här rutan om du vill skriva på dubbla rader i området med de markerade tecknen.  
Inneslutande tecken  
Här definierar du inledande tecken och sluttecken för området med dubbla rader.  
Om du väljer Fler tecken... öppnas dialogrutan Specialtecken där du kan välja bland fler tecken.  
Inledande tecken  
Välj ett inledande tecken för området med dubbla rader.  
Sluttecken  
Välj ett sluttecken för området med dubbla rader.  
Asiatisk typografi  
Här kan du göra några asiatiska typografiska specialinställningar för en cell ett stycke.  
I HTML-dokument går det inte att välja de här alternativen.  
Radbrytning  
Här väljer du de asiatiska typografiska alternativen för radbrytning.  
Använd lista med förbjudna tecken i början och slutet av rader  
Markera den här rutan om du vill att tecknen som inte är tillåtna i början och slutet av rader ska brytas.  
Du matar in listan under Verktyg - Alternativ - Språkinställningar - Asiatisk layout.  
Tillåt hängande interpunktion  
Markera den här rutan om du vill att skiljetecknen som motsvarar komma och punkt inte ska brytas till nästa rad, utan finnas kvar på samma rad - eventuellt även ute i högermarginalen.  
Använd avstånd mellan asiatisk, latinsk och komplex text  
Markera den här rutan om du vill att ett avstånd infogas automatiskt mellan asiatisk, latinsk och komplex text.  
Stycke  
Den här funktionen använder du när du ska redigera styckeegenskaper.  
Om du vill ändra alla stycken av samma typ måste du ändra i den aktuella styckeformatmallen.  
Om Du öppnar den nästan identiska dialogrutan Styckeformatmall via snabbmenyn eller Stylist kommer Du till ytterligare flikar med extra inställningsmöjligheter för textattribut.  
Om Du har öppnat Stylist framhävs det aktuella styckeformatet i Stylist-fönstret.  
Indrag och avstånd  
Här kan du ställa in indrag, avstånd och radavstånd för ett stycke.  
I förhandsvisningen ser du hur ändringarna påverkar utseendet.  
Du kan välja olika måttenheter.  
Indrag  
I området Indrag ställer Du in hur långt texten ska dras in från den vänstra kanten av sidan av textramen av textramen till höger eller från den högra kanten till vänster.  
Du kan definiera ett separat indrag för den första raden.  
Om Du anger ett positivt värde för det vänstra indraget kan Du ändå ange ett negativt värde för den första raden (hängande indrag) eftersom värdet för den första raden hänför sig till värdet Från vänster.  
Från vänster  
I det här rotationsfältet ställer du in styckets avstånd från sidans vänstermarginal.  
Då överskrids vänstermarginalen som har ställts in under Format - Sida - Sida.  
I det här rotationsfältet anger du styckets avstånd från textramens vänstra kant.  
För den första raden är detta avståndet mellan punktuppställningstecknet och textramen om inget annat indrag anges för första raden.  
I det här rotationsfältet anger du styckets avstånd från textramens vänstra kant.  
För den första raden är detta avståndet mellan punktuppställningstecknet och textramen om inget annat indrag anges för första raden.  
Första raden  
Här ställer du in hur långt den första raden ska dras in i förhållande till styckets övriga rader (som ställs in med Från vänster) eller (vid negativt värde) hur långt den ska dras ut.  
Om det aktuella stycket innehåller en numrering / punktuppställning bestäms värdet för den första radens indrag av numreringen och inte av stycket.  
Indraget av första raden för numrerade stycken ställer du in i dialogrutan Numrering / punktuppställning under fliken Position under Avstånd till text.  
Automatiskt  
Markera den här rutan om du vill ha automatiskt indrag.  
Hur mycket den första raden dras in beror då på vilken teckenstorlek och vilket radavstånd som används.  
Inställningen i rotationsfältet Första raden ignoreras.  
Från höger  
Här ställer du in hur långt texten ska dras in från högermarginalen på sidan.  
Då överskrids högermarginalen som är inställd under Format - Sida - Sida.  
Här ställer du in hur långt texten ska dras in från textramens högra kant.  
Här ställer du in hur långt texten ska dras in från textramens högra kant.  
Du kan också ställa in indragen med hjälp av musen.  
Välj då Linjal på menyn Visa.  
Avstånd  
I området Avstånd ställer Du in hur mycket fritt område det ska vara över eller under stycket.  
Det första stycket överst på sidan placeras alltid utan det övre avståndet och det sista stycket underst på sidan utan det undre avståndet.  
Om Du har definierat ett övre respektive ett undre styckeavstånd för två stycken som följer på varandra kommer det största avståndet att gälla såvida Du inte har ställt in något annat under Verktyg - Alternativ - Textdokument - Övrigt.  
Överkant  
I rotationsfältet Överkant ställer Du in hur mycket fritt utrymme (i cm, tum eller annan enhet) det ska finnas över stycket.  
Underkant  
I rotationsfältet Underkant ställer Du in hur mycket fritt utrymme (i cm, tum eller annan enhet) det ska finnas under stycket.  
Radavstånd  
I det här området bestämmer du radavståndet för det aktuella stycket eller för alla markerade stycken.  
Alternativen Enkelt, 1,5 rader eller Dubbelt finns också i undermenyerna till snabbmenyn för det aktuella stycket. De kan också aktiveras med hjälp av ikonerna i objektlisten  
Enkelt  
Med det här alternativet återgår du till enkelt radavstånd.  
Här finns inget extra avstånd mellan raderna.  
Du kan också återgå till enkelt radavstånd med tangentkombinationen Ctrl+1.  
1,5 rader  
Med det här alternativet aktiverar du 1,5-radavståndet.  
Här finns en halv rads extra avstånd mellan raderna.  
Du kan också aktivera det 1,5-radiga radavståndet med hjälp av kortkommandot Ctrl+5.  
Dubbelt  
Med detta alternativ aktiverar Du dubbelt radavstånd.  
Här finns en hel rads extra avstånd mellan raderna.  
Du kan också aktivera det dubbla radavståndet med hjälp av kortkommandot Ctrl+2.  
Proportionellt  
När du väljer det här alternativet aktiveras rotationsfältet med, i vilket Du anger avståndet mellan raderna (100% motsvarar Enkelt).  
Minst  
När du väljer det här alternativet, anger du ett minimiavstånd i rotationsfältet med.  
Eget radavstånd  
I rotationsfältet med anger du ett avstånd som alltid ska läggas till (avstånd mellan underkanten för en rad och överkanten för nästa rad).  
Fast  
Välj ett fast radavstånd i rotationsfältet med.  
Du måste ange minst 0,25 cm.  
Om raderna överlappar vararandra kommer tecknen att kapas.  
med  
I detta rotationsfält anger Du radavståndet som ett procentuellt värde eller absolut värde i cm, beroende på vilken inställning du har valt.  
Om du använder olika teckenstorlekar inom ett stycke anpassar %PRODUCTNAME radavståndet automatiskt till den största teckenstorleken.  
Om du hellre vill ha samma avstånd för alla rader kan du ange ett värde för alternativet Minst som är tillräckligt stort för den största teckenstorleken som används.  
Register  
I det här området kan du ange att Register ska användas som direkt formatering för de markerade styckena eller styckeformatmallen, förutsatt att du har aktiverat det under Format - Sida - Sida.  
Ta hänsyn till  
Markera den här rutan om du vill att register ska användas för styckeformatmallen resp. för alla markerade stycken.  
Tabulator  
Här anger du med numerisk precision tabbarnas placering för stycket.  
Du kan också definiera utfyllnadstecken som ska stå framför tabben på raden.  
Men det kan du bara göra med musen och därför kan du inte göra inställningarna med numerisk precision.  
Position  
I denna ruta anger Du också nya tabbar.  
Dessa är inställda med 2 cm avstånd.  
När Du definierar den första egna tabbplaceringen raderas de standardtabbar som står till vänster.  
I textfältet anger du en tabbplacering i siffror.  
Ange en tabb om 2 cm som 2 eller 2 cm eller 2cm.  
Om du vill använda måttet tum kan du ange 1 tum som 1 ".  
Tryck inte på Retur efter inmatningen - då stängs dialogrutan.  
Klicka i stället på Ny.  
Därefter kan du ange fler tabbar eller ändra typ och utfyllnadstecken för den markerade tabben.  
I den här listrutan finns alla hittills definierade tabbar.  
Du kan markera dem var och en och därefter ändra deras typ och utfyllnadstecken eller radera dem.  
Typ  
I det här området ändrar du typen för den tabb som du har markerat i området Position.  
Vänster  
En vänstertabb är förinställd.  
Text och tal vänsterjusteras till detta läge.  
Höger  
Text och tal högerjusteras till en högertabb.  
Centrera  
Text och tal centreras till en centrerad tabb.  
Decimal  
En decimaltabb vänsterjusterar text medan tal justeras vid det inställda decimaltecknet.  
I den svenska versionen av %PRODUCTNAME är det ett komma.  
Om du anger ett tal (eller ett ord) med decimalkomma justeras talet så att kommat står vid tabulatorn.  
Skiljetecknet för decimalerna styrs av de nationella inställningarna i kontrollpanelen där du kan ändra dem.  
Tecken  
Här anger du det tecken som decimaltabbarna ska justeras vid.  
Det är ett komma i den svenska versionen av %PRODUCTNAME.  
Men du kan även använda andra tecken, t.ex. gradtecken.  
Detta beror på operativsystemet och den teckenuppsättning som används.  
Utfyllnadstecken  
Här väljer Du de utfyllnadstecken som ska infogas före den tabb som Du har markerat under Placering, såvida det inte finns någon annan text där.  
Inga  
Här infogas inga utfyllnadstecken.  
.......  
Här infogas punkter som utfyllnadstecken.  
----- -  
Här infogas bindestreck som utfyllnadstecken.  
______  
Här infogas understrykningstecken som utfyllnadstecken.  
Tecken  
Här används tecken som Du själv har definierat som utfyllnadstecken.  
Tecken  
Ange önskat utfyllnadstecken här.  
Nytt  
När Du har angett ett nytt värde i textfältet Placering aktiveras knappen Ny.  
Genom att klicka på Ny överför Du den nya tabben, inklusive inställningarna för typ och utfyllnadstecken, till listrutan Placering.  
Radera alla  
Med denna knapp raderar Du alla tabbar som finns i listrutan Placering.  
Därefter gäller standardtabbarna, dvs (vänsterjustering, inga utfyllnadstecken, med avståndet 2 cm).  
Inramning  
Under fliken Inramning kan du definiera en inramning för de markerade cellerna det markerade objektet eller det aktuella stycket.  
Du kan tilldela inramningen på alla fyra sidor samma eller olika linjestilar och linjefärger.  
I tabeller kan du även definiera stilen för de inre linjerna.  
Det markerade objektet kan även förses med skuggning.  
Du kan definiera inramningar för sidor, ramar, grafikobjekt, %PRODUCTNAME -tabeller, stycken och integrerade objekt.  
För tabeller i textdokument placerar du markören i tabellen utan att markera något.  
Om du ändrar inramningen nu gäller det för hela tabellen.  
Om du bara vill ha inramning för den aktuella cellen ska du markera den först. (Du måste först markera två celler bredvid varandra med muspekaren och sedan dra tillbaka markeringen till den berörda cellen.)  
Linjeplacering  
Välj en av de fördefinierade inramningarna eller definiera olika linjestilar och linjefärger för varje element i inramningen interaktivt.  
I det övre området kan du snabbt välja de mest använda inramningstyperna.  
Den valda inramningen visas i den grafiska visningen i det undre området där du kan fortsätta att redigera den.  
Du kan även lägga in en inramning genom att använda ikonen Inramning på objektlisten.  
Då öppnas en utrullningslist där du kan välja bland fördefinierade inramningar.  
Inramningen förhandsvisas i det undre fältet.  
De fyra ytterkanterna markeras med små vinklar i det här fältet.  
Om du vill redigera en ytterkant klickar du på motsvarande ställe mellan de små vinklarna.  
De representerar de horisontella och vertikala linjerna mellan cellerna.  
Om du klickar exakt mitt i förhandsvisningen av ramen kan du markera både de inre horisontella och vertikala linjerna samtidigt.  
De element i inramningen som markerats på detta sätt framhävs med svarta trianglar.  
Om du nu väljer en linjestil eller färg gäller ändringen för de markerade elementen i inramningen.  
Om du väljer en tom linje i förhandsvisningen, d.v.s. "ingen linje" visas i stället för "linje "eller "grå linje", så betyder det att den motsvarande delen i inramningen raderas.  
Under fliken Inramning kan du växla cykliskt mellan tre olika tillstånd genom att klicka på ett element upprepade gånger:  
Elementet visas som linje  
Om du avslutar med OK ges elementet den här formateringen.  
Elementet visas som tjock, grå linje  
Om du avslutar med OK ändras inte elementet.  
Elementet visas inte  
Om du avslutar med OK raderas elementet.  
Linje  
I det här området bestämmer du typ och färg för de element i inramningen som är markerade med små trekanter i fältet Ram.  
Den linjestil och linjefärg som du väljer här gäller för de element i inramningen som är markerade i fältet Ram.  
I den övre listrutan finns fördefinierade solida linjer och dubbellinjer med olika linjebredder.  
Välj linjebredd och linjetyp här.  
Alternativet "Ingen" innebär att linjen i det markerade inramningselementet tas bort.  
Om du vill ändra linjestil klickar du på ikonen Linjestil.  
Du väljer linjefärg i kombinationsfältet Färg.  
Svart är förinställd.  
Den valda färgen tilldelas alla markerade inramningslinjer.  
Om du vill ändra linjefärg kan du även klicka på ikonen Ramlinjefärg.  
Avstånd till innehåll  
I det här området definierar du avstånden mellan inramningen och innehållet.  
Om du ökar avstånden leder det till att den tillgängliga platsen för innehållet minskar.  
Det här området visas bara under Format - Sida, men inte under Format - Cell.  
Vänster  
Här anger du textinnehållets avstånd från den vänstra inramningen.  
Höger  
Här anger du textinnehållets avstånd från den högra inramningen.  
Uppe  
Här anger du textinnehållets avstånd från den övre inramningen.  
Nere  
Här anger du textinnehållets avstånd från den nedre inramningen.  
Synkronisera  
Om du markerar den här rutan, får alla fyra avstånden samma värde nästa gång du ändrar ett avstånd.  
Skuggning  
Du kan förse inramningen med en skuggning, som läggs bakom inramningen på två bredvidliggande sidor.  
Det sker oavsett om själva inramningen syns.  
Om grafikobjektet eller objektet i dokumentet är förankrat i en textram så kan grafikobjektet eller objektet inte sträcka sig utanför textramens kant.  
Detta gäller inklusive skuggning.  
Om ett objekt, som fyller hela textramen utan skuggning, förses med skuggning, trycks objektet ihop så pass mycket att även skuggningen får plats i textramen.  
Position  
Välj en av de fördefinierade skuggningsvarianterna här.  
Den valda skuggningen visas under Ram.  
Distans  
Ange önskad distans för skuggan här.  
Färg  
Välj önskad skuggfärg här.  
Bakgrund  
Här definierar du bakgrundsfärg eller väljer en bakgrundsbild.  
Du kan definiera de här egenskaperna för stycken, sidor, sidhuvuden och sidfötter, textramar, tabellceller och tabeller, områden och förteckningar i det aktuella stycket eller i markerade stycken.  
Definiera bakgrundsfärg för celler och dessutom en bakgrundsbild för sidformatmallen.  
som  
Här anger Du om det är en bakgrundsfärg eller en bakgrundsbild som ska redigeras.  
Om Du väljer Grafik, kan Du ange en viss bild som bakgrund.  
Om Du öppnar den här dialogrutan med menykommandot Format - Tecken... eller Format - Cell... eller Format - Objekt... kan Du inte använda kombinationsfältet Som.  
Den dialogruta som motsvarar valet Som Färg öppnas.  
Om du har valt färgen:  
Bakgrundsfärg  
Välj en färg som bakgrundsfärg eller klicka på "Ingen fyllning".  
Nedanför färgrutorna visas namnet på den aktuella bakgrundsfärgen.  
Område  
Här anger Du för vilket område den valda bakgrundsfärgen ska gälla.  
Om det är fråga om en bakgrundsfärg för en styckeformatmall kan Du här välja om färgen ska gälla stycket eller de markerade tecknen.  
Om det är fråga om en tabell anger Du om färgen ska gälla den aktuella cellen, den aktuella raden eller hela tabellen.  
Det här kombinationsfältet visas bara om bakgrundsfärgen gäller en tabell eller en styckeformatmall.  
Om Du har valt Som Grafik:  
Fil  
Du kan också söka i filer och skapa länkar.  
Fil:  
Här får Du information om länkar till grafikobjektet.  
Länka  
Här kan Du länka det markerade grafikobjektet till dokumentet.  
Förhandsvisning  
Markera den här rutan om du vill titta på det valda grafikobjektet i förhandsvisningen innan du integrerar det i dokumentet  
Välj ut...  
Om du trycker på den här kommandoknappen kommer du till dialogrutan Sök grafik.  
Den är uppbyggd på ungefär samma sätt som dialogrutan Infoga grafik.  
Typ  
Här definierar du visningstyp för bakgrundsgrafiken.  
Position  
När du har valt Position, definierar du grafikens position på sidan i det tillhörande förhandsvisningsfältet.  
Yta  
Om du väljer alternativet Yta, infogas grafikobjektet en gång bakom det objekt för vilket du har definierat bakgrunden.  
Om Du väljer det här alternativet, inpassas den markerade bilden i ett exemplar på ytan och i förekommande fall förvriden.  
Sida vid sida  
Om Du väljer alternativknappen Sida vid sida, upprepas bilden i ett rutmönster bakom objektet (tabellen, textramen, sidan osv) och varje förekomst infogas i originalstorlek.  
Här väljer du en färg från färgpaletten.  
Justering  
Här kan du ställa in justeringen för ett stycke.  
Justering  
I detta område anger Du om stycket ska vänster - eller högerjusteras, centreras eller marginaljusteras.  
Dessa alternativ finns också i det aktuella styckets snabbmeny.  
Du kan också använda ikonerna på objektlisten.  
Vänster  
Med detta alternativ vänsterjusterar du stycket.  
Höger  
Med det här alternativet högerjusterar du stycket.  
Centrerat  
Med det här alternativet centrerar du stycket.  
Marginaljustering  
Med det här alternativet marginaljusterar du stycket.  
Vid marginaljustering dras alla rader i stycket (förutom sista raden) ut till samma bredd.  
På så sätt undviker du att marginalen blir ojämn.  
Det här alternativet används ofta när en sida innehåller flera spalter.  
Sista raden  
Här definierar Du hur den sista raden i marginaljusteringen ska formateras.  
Du kan välja mellan Vänster, Centrerad och Marginaljusterad.  
Expandera enstaka ord  
Här kan Du välja att dra ut ett ord, som är det enda som står på den sista raden men som hör till ett stycke som marginaljusterats, över hela raden.  
Detta görs genom att avståndet mellan bokstäverna förstoras.  
Detta fungerar dock endast om Du valt Marginaljusterad i rutan Sista raden.  
Ersätt då blankstegen i raden med skyddade blanksteg genom att trycka på Kommando Ctrl och mellanslag.  
Vertikal textjustering  
Välj här förinställningarna för den vertikala justeringen av texttecken på textraden.  
Du kan välja bland Automatiskt, Baslinje, Uppe, Centrerat och Nere.  
Du ser t.ex. effekten om du formaterar några tecken i ett stycke i en betydligt större teckenstorlek än de andra.  
Beskära  
Här kan du beskära visningen av ett grafikobjekt samt definiera dess storlek och skala.  
Själva grafikobjektet förändras inte; de här inställningarna påverkar bara den aktuella visningen av objektet.  
Beskär  
I det här området ändrar du visningen av grafikobjektet - positiva värden förstorar marginalen mellan ram och objekt medan negativa värden beskär grafikobjektet.  
Om du anger negativa värden ser du en ram i förhandsvisningsfönstret som visar vilket område av grafikobjektet som finns kvar och vad som tas bort.  
Bibehåll skalning  
Om Du vill att proportionerna mellan grafikobjektets sidor ska behållas efter beskärningen - för att undvika att det förvrängs - markerar Du det här alternativfältet.  
Med det här alternativet innebär en beskärning bara att storleken ändras.  
Grafikobjektets skala ändras inte.  
Bibehåll bildstorlek  
Klicka här om grafikobjektets ursprungliga storlek ska behållas efter beskärningen.  
Med det här alternativet innebär en beskärning bara att skalan ändras.  
Grafikobjektets storlek ändras inte.  
Vänster  
Här definierar du med hur mycket den vänstra sidan av det markerade grafikobjektet ska ändras.  
Höger  
Här bestämmer du med hur mycket den högra sidan av det markerade grafikobjektet ska ändras.  
Uppe  
Här anger du med hur mycket den övre kanten av det markerade grafikobjektet ska ändras.  
Nere  
Här definierar du med hur mycket underkanten av det markerade grafikobjektet ska ändras.  
Skalning  
I det här området kan du ändra grafikobjektets bredd och höjd.  
Om du gör en ändring i området Skala sker en proportionell anpassning i området Storlek.  
Bredd  
Här definierar du det aktuella grafikobjektets bredd.  
Inmatningen görs i procent.  
Höjd  
I det här rotationsfältet definierar du grafikobjektets höjd.  
Inmatningen görs i procent.  
Bildstorlek  
I det här området kan du ändra grafikobjektets bredd och höjd.  
Om du gör en ändring i området Storlek sker en proportionell anpassning i området Skala.  
Bredd  
I det här rotationsfältet definierar du grafikobjektets bredd.  
Höjd  
I det här rotationsfältet definierar du grafikobjektets höjd.  
Originalstorlek  
Om Du klickar på den här kommandoknappen återkallas ändringarna i områdena Skala och Storlek, och grafikobjektets originalstorlek återställs.  
Administrera  
Under den här fliken administrerar du en formatmall.  
Om du vill göra ett dokument till dokumentmall, använder du kommandot Arkiv - Dokumentmall - Spara.  
Om du vill överföra formatmallar från ett visst dokument till det aktuella dokumentet, använder du kommandot Format - Mallar - Ladda.  
Om du rent allmänt vill kopiera eller flytta formatmallar från ett dokument till andra mallkategorier eller dokument, använder du kommandot Format - Mallar - Katalog.  
Namn  
Här visas namnet på formatmallen.  
Om du skapar en ny formatmall, anger du dess namn här.  
Det kan bestå av upp till 256 kombinerade bokstäver, siffror och specialtecken.  
Om det redan finns en mall med det namn som du anger, visas ett meddelande om detta.  
Det går alltså inte att välja textfältet i det här fallet.  
Det är bara användardefinierade mallar som kan döpas om.  
Automatisk uppdatering  
Om du markerar den här rutan uppdateras formatmallen automatiskt när ett objekt ändras, precis som när du klickar på Uppdatera mall i Stylist.  
Nästa formatmall  
Klicka i kombinationsfältet och välj namnet på önskad formatmall.  
Först är det aktuella mallnamnet markerat.  
När det gäller styckeformatmallar infogas bara nästa formatmall automatiskt när du trycker på returtangenten.  
När det gäller formatering i efterhand måste du göra tilldelningen för hand.  
För sidformatmallar verkställs den angivna formateringen enligt Nästa formatmall automatiskt vid sidbrytningen.  
Den här funktionen är bara tillgänglig för stycke - och sidformatmallar.  
Länkad med  
Klicka i fältet och välj den mall med vilken den aktuella mallen ska vara länkad.  
Formaten i den länkade mallen används som bas för formaten i den aktuella mallen.  
Den här funktionen är bara tillgänglig för stycke-, tecken - och ramformatmallar.  
Kategori  
Här visas den mallkategori som den aktuella mallen tillhör.  
När du skapar en ny formatmall, klickar du i det här fältet och väljer mallkategori.  
För användardefinierade mallar är det lämpligt att välja posten Användardefinierade formatmallar, så att du undviker förväxlingar med de mallar som följer med programmet.  
Det går alltså inte att aktivera kombinationsfältet i det här fallet.  
Innehåller  
Här visas skillnaderna mellan formatmallen och inställningarna från den överordnade formatmallen.  
För några typer av formatmallar räknas alla egenskaper upp här.  
Sida  
Här definierar du marginaler, olika layouter för flersidiga dokument, numrering samt pappersformat.  
Du göra olika standardinställningar, t.ex. för det pappersformat som ska användas, pappersorientering, utskriftsområde och sidlayout.  
Du kan använda olika måttenheter.  
Pappersformat  
Här finns ett urval vanliga pappersformat.  
Om du definierar ett pappersformat här, visas automatiskt tillhörande mått i rotationsfälten Bredd och Höjd.  
Format  
Välj ett fördefinierat format i listrutan Format för utskrift på papper eller bildskärm.  
Den här funktionen är praktisk för bildskärmspresentationer och HTML-sidor.  
Här kan du ange en pappersbredd som avviker från förinställningen.  
Höjd  
Här kan du ange en pappershöjd som avviker från förinställningen.  
Stående  
Välj det här alternativet om dokumentet ska skrivas ut i stående format (höjdformat).  
Liggande  
Välj det här alternativet om dokumentet ska skrivas ut i liggande format (landscape).  
Pappersmatning  
Om din skrivare har flera fack för pappersinmatning, kan du definiera vilket av dem som ska användas här.  
Om papperstypen ska bytas efter första sidan måste du ange vilka fack som ska användas.  
Välj skrivarfack för första arket i dialogrutan Skriv ut och för andra och följande ark i dialogrutan Format - Sida.  
Detta förutsätter att du för sidan 2 och följande sidor har definierat en annan sidformatmall än för sidan 1.  
Sidmarginaler  
Du kan definiera avståndet mellan textytan och pappersarkets kant.  
Standardinställningen är 2 cm.  
De här värdena är i samtliga fall större än minimimåttet för alla gängse skrivarmodeller och garanterar därmed att ingen del av dokumentet faller bort vid utskriften.  
Du kan ändra marginalmåtten i rotationsfälten.  
Här kan du även ange olika måttenheter, och måtten räknas då automatiskt om.  
Vänster / Inre  
I det här anger rotationsfältet kan du definiera bredden på vänster respektive inre marginal.  
Om du har valt sidlayouten Spegelvänt, heter det här rotationsfältet Inre och anger den inre marginalen vid dubbelsidig utskrift.  
Höger / Yttre  
Här kan du definiera bredden på höger respektive yttre marginal.  
Om du har valt sidlayouten Spegelvänt, heter det här rotationsfältet Yttre och anger den yttre marginalen vid dubbelsidig utskrift.  
Uppe  
Här bestämmer du den övre marginalens storlek.  
Nere  
Här bestämmer du den nedre marginalens storlek.  
Om du ställer in och bekräftar (med OK) marginaler som är sådana att en del av sidan faller utanför det utskrivbara området, blir du upplyst om detta i en dialogruta där du även blir uppmanad att bekräfta inställningarna igen.  
Du kan ångra inställningarna med kommandoknappen Nej.  
I så fall ersätts de ogiltiga värdena automatiskt med giltiga, som läggs så nära dem som du har angett som möjligt.  
Då visas det maximala respektive minimala marginalmåttet.  
Layoutinställningar  
När du väljer sidlayout bestämmer du hur mycket layouten ska omfatta.  
Sidlayout  
I det här kombinationsfältet definierar du på vilka sidor i dokumentet som inställningarna ska gälla.  
Höger och vänster  
Inställningarna kommer att användas på alla sidor i dokumentet.  
Spegelvänt  
Den här sidlayouten är avsedd för dokument med dubbelsidig utskrift, där arken ska häftas eller bindas in.  
Bara höger  
Inställningarna används bara på högersidor.  
Dokumentets första sida är automatiskt en högersida.  
Bara höger  
Inställningarna används bara på vänstersidor.  
Register  
Här aktiverar och inaktiverar du Register.  
Det här området finns bara i formatdialogrutan för stycken och sidor, däremot inte för ramar med flera kolumner.  
Aktivera  
Om du vill aktivera register för alla sidor i den här mallen markerar du den här rutan.  
Referensstyckeformatmallen bestämmer radhöjden för rastret.  
Referensstyckeformatmall  
Välj den styckeformatmall i listrutan som ska vara standardmall.  
I alla stycken där register är aktiverat justeras alla rader med sina baslinjer så som baslinjerna är justerade i ett stycke, som är formaterat med referensstyckeformatmallen.  
Tabelljustering  
I det här området definierar du justering av cellinnehållet.  
Horisontellt  
Markera den här rutan om du vill ha en horisontellt centrerad orientering.  
Vertikalt  
Markera den här rutan om du vill ha en vertikalt centrerad orientering.  
Layoutinställningar  
Format  
I det här kombinationsfältet väljer du typ av sidnumrering.  
Anpassa till storlek  
Här kan du ange om du även vill behålla teckningselementens placering om pappersformatet ändras.  
Om den här rutan är markerad, placeras alla objekt innanför marginalerna om om sidstorleken ändras så att sidlayouten inte ändras.  
Speciellt anpassas placeringen, storleken och, i fråga om presentationsobjekt på sidformatmallen (masterpage), mallens teckenstorlek till den nya layouten.  
På detta sätt kan du t.ex. avbilda sidlayouten i en mall på olika sidformat.  
Sidhuvud  
Här lägger du in ett sidhuvud för dokumentet och definierar dess egenskaper.  
Sidhuvuden är områden som är åtskilda från arbetsområdet, är fast förankrade och upprepas överst på varje sida.  
Oberoende av arbetsområdet kan de förses med en bakgrund och även ramas in.  
Du kan använda olika måttenheter.  
För att kunna foga in och ta bort ett sidhuvud på alla sidor som försetts med en viss sidformatmall kan Du även välja kommandot Infoga - Sidhuvud.  
Ramar i sidhuvuden och sidfötter som är bundna till stycken får sträcka sig över satsytan, både till vänster och till höger.  
Om du vill ta med grafikobjekt och andra objekt i huvudet på varje utskriven sida fogar du in dessa på tabellens första rad (t.ex. i cellen A1).  
Raden skrivs ut automatiskt på varje sida i dokumentet.  
Med tangentkombinationen Ctrl+PageUp växlar du mellan text och sidhuvud.  
Med kortkommandona Ctrl+PageUp och Ctrl+Page Down växlar Du fram och tillbaka mellan sidhuvud och sidfot.  
Sidhuvud  
Här kan olika inställningar för sidhuvudet göras, t ex sidhuvudets höjd och radavstånd.  
Sidhuvud på  
Om du vill förse dokumentet med ett sidhuvud markerar du den här rutan.  
Avstånd  
I det här rotationsfältet anger du önskat avstånd till texten.  
Höjd  
I detta rotationsfält anges den önskade höjden på sidhuvudet.  
Anpassa höjd dynamiskt  
Markera den här rutan om du vill att sidhuvudets höjd ska anpassas dynamiskt till textmängden och den använda teckenstorleken i sidhuvudet.  
Vänstermarginal  
Här anges avståndet mellan sidhuvudets vänsterkant och papperets vänsterkant.  
Högermarginal  
Här anges avståndet mellan sidhuvudets högerkant och papperets högerkant.  
Samma innehåll höger / vänster  
Avmarkera den här rutan om du behöver olika sidhuvuden på höger och vänster sida för dokument med dubbelsidigt tryck.  
Om du inte har gjort någon markering är sidhuvudena för vänster och höger sida olika.  
Om du klickar på kommandoknappen Redigera kan du definiera innehållet för höger - och vänstersidor separat.  
Fler...  
Under Fler kan Du definiera en ram eller annan bakgrund bakom sidhuvudet.  
Du kommer till dialogrutan Inramning / Bakgrund med flikarna Inramning och Bakgrund.  
Redigera...  
Med denna kommandoknapp öppnar Du en dialogruta för att redigera sidhuvud eller sidfot.  
Sidfot  
Här väljer du en sidfot och definierar deras placering.  
En sidfot är ett område som är åtskilt från arbetsområdet, är fast förankrat och upprepas längst ner på varje sida.  
Den kan förses med en annan bakgrund än arbetsområdet och ramas in av en linje.  
Du kan använda olika måttenheter.  
Om Du vill infoga eller ta bort en sidfot på alla sidor som använder en bestämd sidformatmall kan Du använda kommandot Infoga - Sidfot.  
Ramar i sidhuvuden och sidfötter som är bundna till stycken kan Du låta sträckas ut över satsytan, både till höger och till vänster.  
Med hjälp av tangenterna Ctrl+Page Down växlar Du mellan texten och sidfoten.  
Med tangenterna Ctrl+Page Up och Ctrl+Page Down växlar Du mellan sidhuvudet och sidfoten om sådana finns.  
Sidfot  
Du kan t ex ställa in sidfotshöjden eller kantavstånden.  
Sidfot på  
Markera den här rutan om du vill förse dina dokument med en sidfot.  
Avstånd  
I detta rotationsfält anger Du det önskade avståndet till brödtexten.  
Höjd  
I detta rotationsfält anger Du önskad höjd för sidfoten.  
Anpassa höjden automatiskt  
Markera den här rutan om du vill att sidfotens höjd ska anpassas dynamiskt till textmängden och den använda teckenstorleken i sidfoten.  
Vänstermarginal  
Här definierar Du det avstånd som sidfotens vänstermarginal ska dras in i förhållande till den vänstra textmarginalen.  
Högermarginal  
Här definierar Du det avstånd som sidfotens högermarginal ska dras in i förhållande till den högra textmarginalen.  
Samma innehåll höger / vänster  
Avmarkera den här rutan om dokument som skrivs ut på båda sidor ska ha olika sidfotstexter på vänster - respektive högersidor.  
Om du inte har markerat den här rutan kommer sidfötterna att vara olika för höger - respektive vänstersidor.  
Genom att klicka på kommandoknappen Redigera definierar du innehållet för höger - respektive vänstersidor separat.  
Tillägg...  
Under Tillägg definierar Du en inramning eller annan bakgrund för sidfoten.  
Dialogrutan Inramning / bakgrund med flikarna Inramning och Bakgrund visas.  
Redigera...  
Med denna knapp kommer Du till dialogrutan Redigera - Sidhuvud och sidfot.  
Bokstäver / tecken  
Med kommandona på den här undermenyn omvandlar du den markerade texten eller ordet under markören.  
Stora bokstäver  
Omvandlar västlig text till stora bokstäver.  
Små bokstäver  
Omvandlar västlig text till små bokstäver.  
Halv bredd  
Omvandlar asiatisk text till halv bredd.  
Normal bredd  
Omvandlar asiatisk text till normal bredd.  
Hiragana  
Omvandlar text till Hiragana.  
Katakana  
Omvandlar asiatisk text till katakana.  
Ruby  
I dialogrutan Ruby matar du in kompletterande text som är tilldelad den markerade texten.  
Ruby är beteckningen för en text som står direkt ovanför eller nedanför en annan text (bastext) och som innehåller en anmärkning eller förklaring av uttalet.  
Markera ett eller flera ord i ett dokument.  
Välj Format - Ruby.  
Ange ruby-texten till varje ord.  
Bastext  
I det här området ser du bastexten som en Ruby-text ska användas för.  
Ruby-text  
Här skriver du respektive ruby-text för bastexten.  
Justering  
Här bestämmer du justeringen.  
Position  
Här väljer du var ruby-texten ska placeras.  
Teckenformatmall för ruby-text  
Välj vilken teckenformatmall du vill använda för ruby-texten.  
Stylist  
Med den här kommandoknappen öppnar du Stylist Stylist.  
Justering (objekt)  
Den här funktionen använder du för att justera objekt.  
De olika justeringsalternativen beror på objekttypen och förankringen.  
Multipel markering påverkar också.  
Exempelvis justeras bara flera markerade teckningselement eller kontrollfält i förhållande till varandra om de är förankrade vid sidan eller stycket och inte om de är förankrade som tecken.  
Med den här ikonen kan du dra upp ett fönster och flytta bort det från listen.  
I fönstret hittar du ikoner för alla de justeringsfunktioner som beskrivs här.  
Vänster  
Flera markerade objekt justeras mot vänstra kanten på det objekt som är placerat längst till vänster.  
Om objektet är förankrat på sidan, i ett stycke, tecken eller ram, vänsterjusteras det i förhållande till referenselementet.  
Vid förankring som tecken är denna funktion inte tillgänglig.  
Referenselementet kan t.ex. vara ett styckeområde eller hela sidan.  
Det definieras under fliken Typ.  
Om flera element är markerade, t.ex. teckningselement eller kontrollfält, justeras de in med sin vänstersida mot den objektsida som är placerad längst till vänster.  
Denna relativa justering sker endast vid multipel markering, inte om respektive element är grupperade.  
Grupperade element fungerar som ett enda objekt vid justering.  
Centrerad  
Flera markerade objekt justeras med mittpunkten på en linje.  
Om objektet är förankrat vid sidan, vid stycket, vid tecknet eller vid ramen justeras det horisontellt centrerat i förhållande till referenselementet.  
Denna funktion är inte tillgänglig för förankring som tecken.  
Om du har markerat flera element, t.ex. teckningselement eller kontrollfält, justeras de horisontellt centrerat i förhållande till varandra så att deras mittpunkter ligger ovanpå varandra.  
Den vertikala positionen påverkas inte.  
Höger  
Flera markerade objekt justeras mot högra kanten på det objekt som är placerat längst till höger.  
Om objektet är förankrat på sidan, i ett stycke, tecken eller ram, högerjusteras det i förhållande till referenselementet.  
Denna funktion finns inte tillgänglig för förankring som tecken.  
Om flera element är markerade, t.ex. teckningselement eller kontrollfält, justeras de in med sin högersidor mot den objektsida som är placerad längst till höger.  
Uppe  
Flera markerade objekt justeras vid den övre kanten på det objekt som står längst till upp.  
Om objektet är förankrat vid sidan, stycket, tecknet eller ramen justeras det i förhållande till referenselementet på så sätt att dess övre kant orienteras efter referenselementets övre kant.  
Detta gäller även om du har valt förankringen "som tecken".  
Men om du väljer baslinjen som referenselement, sätts den undre kanten på objektet på linjen där alla tecken på raden står (baslinje).  
Referenselementet kan t.ex. vara ett textområde.  
Det definieras under fliken Typ.  
Om flera element är markerade, t.ex. teckningselement eller kontrollfält, justeras alla med sina övre sidor vid den objektsida som är placerad högst upp.  
Centrerat  
Om flera objekt är markerade justeras de med sina mittpunkter på en vertikal linje.  
Om objektet är förankrat till sidan, till ett stycke, till ett tecken, som tecken eller till en ram, centreras det vertikalt i förhållande till referenselementet.  
Om flera element är markerade, t.ex. teckningselement eller kontrollfält, justeras de vertikalt centrerat i förhållande till varandra på så sätt att deras mittpunkter ligger på samma höjd.  
Den horisontala placeringen påverkas inte.  
Underst  
Flera markerade objekt justeras in mot underkanten på det objekt som är placerat underst.  
Den undre kanten på objektet orienterar sig efter den undre kanten på referenselementet.  
Detta gäller även vid förankring "som tecken".  
Men om du väljer baslinjen som referenselement sätts objektets övre kant på den linje där alla tecken på raden står (baslinje).  
Om flera element är markerade, t.ex. teckningselement eller kontrollfält, justeras de med sina undre sidor mot den objektsida som är placerad längst ned.  
Justering (textobjekt)  
Det här kommandot visar alla möjligheter att justera textobjekt.  
Info: du får ett textobjekt om du dubbelklickar på en teckning som du har skapat med ritfunktionerna.  
Vänster  
Med kommandot Vänster eller ikonen Vänsterjusterat gör du det aktuella stycket vänsterjusterat.  
Om flera stycken är markerade, gäller kommandot för alla markerade stycken.  
Höger  
Med kommandot Höger eller ikonen Högerjusterat högerställer du det aktuella stycket.  
Om flera stycken är markerade gäller kommandot samtliga markerade stycken.  
Centrerat  
Med detta kommando centreras texten i det aktuella stycket.  
Om flera stycken är markerade gäller kommandot för samtliga markerade stycken.  
Marginaljustering  
Med det här kommandot dras alla rader i det aktuella stycket ut till samma längd.  
Den sista raden behandlas för sig (ställ in detta under Format - Stycke - Justering).  
Om flera stycken är markerade, gäller kommandot för alla.  
Teckensnitt  
Med detta kommando ser du alla teckensnitt som kan väljas när du har markerat ett textobjekt.  
Info: du får ett textobjekt om du dubbelklickar på en teckning som du har skapat med ritfunktionerna.  
Storlek  
Det här kommandot visar alla teckenstorlekar som kan väljas för ett aktiverat textobjekt.  
Info: du får ett textobjekt om du dubbelklickar på en teckning som du har skapat med ritfunktionerna.  
Stil  
Med det här kommandot visas de viktigaste möjligheterna att ge textobjekt effekter och tilldela dem en teckenstil.  
Info: du får ett textobjekt om du dubbelklickar på en teckning som du har skapat med ritfunktionerna.  
Med den här funktionen kan du snabbt nå de viktigaste kommandona från fliken Format - Tecken - Teckensnitt och Format - Tecken - Teckeneffekt.  
Om markören befinner sig i ett ord, formateras hela ordet om.  
Om bara ett eller flera tecken är markerade, gäller kommandot just dem.  
Om ingenting är markerat, och markören inte står i något ord, gäller den valda stilen de tecknen som skrivs in därefter.  
Fet  
Med det här kommandot formaterar du den markerade texten, eller ordet som markören står i, med fetstil.  
Om textmarkören inte står i ett ord formateras all den text som du skriver när du har tryckt på ikonen Fet med fetstil tills du trycker på ikonen igen eller flyttar markören.  
Kursiv  
Med detta kommando kursiverar du den markerade texten eller det ord som markören står i.  
Om textmarkören inte står i ett ord kursiveras all den text som du skriver när du har tryckt på ikonen Kursiv tills du trycker på ikonen igen eller flyttar markören.  
Understruken  
Med kommandot Understruken eller ikonen Understruken stryker du under den markerade texten eller det ord i vilken markören befinner sig.  
Om textmarkören inte står i ett ord stryks den text under som du skriver när du har klickat på ikonen Understruken tills du klickar på ikonen igen eller flyttar markören.  
Med kommandot Dubbelt understruken stryks tecknen under dubbelt.  
Genomstruken  
Med det här kommandot stryker du igenom den markerade texten eller det ord där markören står.  
Skuggad  
Med detta kommando visas den markerade texten eller det ord, i vilket markören står, med skuggning.  
Kontur  
Via detta kommando förses den markerade texten, eller det ord där markören står, med en kontur.  
Upphöjt  
Med det här kommandot gör du den markerade texten, eller det ord där markören står, upphöjd.  
Nedsänkt  
Med detta kommando sänks den markerade texten, eller det ord där markören står, ned.  
Radavstånd  
Det här kommandot visar de viktigaste inställningarna som är möjliga för radavstånd i textobjekt.  
Info: du får ett textobjekt om du dubbelklickar på en teckning som du har skapat med ritfunktionerna.  
Med den här funktionen kan du snabbt nå de viktigaste radavstånden under fliken Format - Stycke - Indrag och Avstånd.  
Enkelt radavstånd  
Med detta kommando ger du det aktuella stycket ett enkelt radavstånd.  
Om flera stycken är markerade gäller kommandot för samtliga markerade stycken.  
1,5 rader  
Med detta kommando ger du det aktuella stycket ett radavstånd på en och en halv rad (1,5).  
Om flera stycken är markerade gäller kommandot för samtliga markerade stycken.  
Dubbelt  
Med det här kommandot definierar du att det aktuella stycket ska ha dubbelt radavstånd.  
Om flera stycken är markerade, gäller kommandot för alla.  
Skapa mall  
Mallens namn  
Här finns ett textfält där Du kan ange namnet på en ny mall och ett fält med en lista som visar alla befintliga mallar.  
Mallens namn  
Skriv ett namn för den nya mallen eller välj ett namn i listrutan nedanför.  
Mallens namn  
I den här rutan visas en lista över befintliga mallar.  
Om Du väljer en mall från listan får Du ett meddelande om att den här mallen redan finns.  
Om Du klickar på Ja skrivs den befintliga mallen över.  
Lägga till AutoFormat  
Namn  
Här anger Du namnet på det nya AutoFormatet.  
Linje  
I dialogrutan Linje ställer du in utseendet för ritade linjer.  
Den här funktionen är bara tillgänglig om du har markerat ett ritat objekt.  
Linje  
Här väljer du en fördefinierad linjestil, färg och bredd.  
Dessutom kan du välja bland fördefinierade linjeslut.  
Linjeegenskaper  
Stil  
Under Format - Linje - Linjestilar kan du definiera egna linjestilar.  
Färg  
I det här kombinationsfältet definierar du linjefärgen.  
Bredd  
Definiera linjebredden här.  
Du kan använda olika måttenheter.  
Transparens  
Här väljer du transparens från 0% (täckande) till 100% (genomskinligt).  
Följande område visas bara under fliken Inramning i dialogrutan Dataserie, om du har valt diagramtypen XY-diagram.  
Symbol  
I det här området kan du välja symboler för datapunkterna i diagrammet.  
Urval...  
På undermenyn kan du välja en symbol.  
Förutom Ingen symbol kan du välja:  
Automatiskt, Från fil, Gallery och Symboler. "Automatiskt" använder de förinställda standardsymbolerna, som också skalas automatiskt. "Från fil... "öppnar dialogrutan Länka, som motsvarar dialogrutan Öppna.  
Där kan du välja en symbol.  
Med "Gallery" väljer du ett av grafikobjekten från Gallery-temat Punkter.  
Under "Symboler" hittar du en lista med förinställda symboler.  
Bredd  
Ställ in symbolbredden här Om du ställer in Automatiskt beräknas värdet ur bredden på förklaringstexten och därför är rotationsfältet inte aktiverat..  
Höjd  
Här ställer du in symbolhöjden.  
Om du har ställt in Automatiskt beräknas värdet ur höjden på förklaringstexten och därför är rotationsfältet inte aktiverat.  
Proportionellt  
Om rutan är markerad ändras även höjden proportionellt om bredden ändras (och tvärtom).  
Linjeslut  
I det högra området kan du välja bland olika linjeslut.  
Under fliken Linjeslut kan du välja fler linjeslut.  
Du kan också definiera egna linjeslutsymboler.  
Stil  
Välj här en av de fördefinierade symbolerna för linjeslut.  
Bredd  
Skriv den önskade bredden på linjeslutsymbolen, eller ställ in önskat värde med pilknapparna.  
Om Du vill upphäva visningen av linjeslutsymbolerna ställer Du in måttet 0,00 cm under Bredd.  
Centrerat  
Med hjälp av kryssrutorna centrerad kan Du placera mitten av linjeslutsymbolen på linjeslutet.  
Linjen förlängs på detta sätt.  
Om denna kryssruta inte är aktiv placeras linjesymbolen på linjen på ett sådant sätt att linjens längd inte förändras.  
Synkronisera slut  
Om Du väljer detta alternativ gäller de inställningar som Du gör för den ena linjeslutsymbolen automatiskt även för den andra symbolen.  
Linjestilar  
Här kan du ändra och själv definiera linjestilar.  
Egenskaper  
Linjestil  
Välj den linjetyp som ska ändras.  
Typ  
Välj kombination här.  
Du kan skapa användardefinierade linjetyper genom att kombinera punkter och streck.  
Heldragna linjer skapar du med en kombination av typerna Bindestreck-Bindestreck.  
Antal  
Ange här det antal punkter eller streck som ska följa på varandra.  
Längd  
Här kan du definiera längden för linjetypen streck.  
Avstånd  
Ange här avståndet mellan de enskilda linjestilarna.  
Anpassa till linjebredd  
Om du markerar den här kryssrutan gäller alla måttangivelser i förhållande till linjebredden.  
Den verkliga linjebredden ställer du in under Format - Linje - Linje.  
Lägg till...  
Om du klickar här öppnas en dialogruta där du kan ange ett namn för en ny linjestil med de aktuella inställningarna.  
Namn  
Skriv namnet här.  
Ändra...  
Om du klickar här öppnas en dialogruta där du kan mata in ett nytt namn för den markerade linjestilen.  
Mata in ett nytt namn eller bekräfta det gamla namnet.  
De aktuella inställningarna används för den markerade linjestilen.  
Ladda linjestilstabell  
Om du klickar på den här ikonen öppnas dialogrutan Öppna där du kan ladda en linjestilstabell.  
Spara linjestilstabell  
Om du klickar på den här ikonen öppnas dialogrutan Spara som där du kan spara en linjestilstabell.  
Linjeslut  
Här definierar eller ändrar du ett linjeslut.  
Administrera linjeslut  
Ange det nya namnet för linjeslutet i det övre textfältet, eller välj ett linjeslut i det nedre kombinationsfältet.  
Linjeslutstil  
I textfältet anger du ett namn för linjeslutet.  
Namn  
I kombinationsfältet väljer du en av de fördefinierade linjesluten.  
Lägg till...  
Här ger du ett teckningselement som du själv har skapat ett namn.  
Du måste först rita teckningselementet med en spets som pekar uppåt, och markera det.  
Ändra...  
Mata in ett annat namn i fältet Namn och klicka på den här kommandoknappen om du vill ändra namnet.  
Ladda linjesluttabell  
Med den här ikonen öppnar du dialogrutan Öppna.  
Spara linjesluttabell  
Med den här ikonen öppnar du dialogrutan Spara som.  
Yta  
Med denna funktion kan du redigera objektytor.  
I dialogrutan kan du definiera ytans egenskaper, färger och gradienter och redigera skrafferingar och bitmappmönster.  
Den här funktionen kan du bara använda när du har markerat ett ritobjekt.  
Yta  
Här bestämmer du om den markerade ytan ska fyllas med en färg, en färggradient, en skraffering eller en bitmap.  
Du kan spara ändrade färger, färggradienter, skrafferingar och bitmap-mönster som användardefinierade filer.  
Fliken heter Bakgrund om du öppnar den i %PRODUCTNAME Impress eller %PRODUCTNAME Draw via Format - Sida.  
Fyllning  
Här väljer du ytfyllningens typ eller färg.  
Först anger du ytstil, och sedan kan du definiera fyllningsmöster och fyllningsfärg för den valda ytstilen i listrutan Ytfyllning.  
Listrutor på objektlisten:  
Ingen  
Du väljer det här alternativet när den aktuella ytfyllningen inte ska visas.  
Om du har gjort ytan osynlig och vill ångra det här attributet, måste du inte bara tilldela den en annan ytstil (t.ex. färg) utan även välja en tillhörande färg.  
I annat fall upphävs inte alternativet Ingen.  
Färg  
Om Du skulle vilja fylla ytan med en färg från den aktuella färgtabellen, klickar Du här.  
Valet gör Du i listrutan Ytfyllning.  
Om du har markerat ett objekt vars färg inte finns med i färgtabellen, visas färgen ändå här.  
I dialogrutan Format - Yta - Färger kan du överta den med Lägg till.  
Färggradient  
Ytan fylls med en färggradient från den aktuella färggradienttabellen.  
Valet gör Du i listrutan Ytfyllning.  
Skraffering  
Ytan fylls med en skraffering från den aktuella skrafferingstabellen.  
Valet gör Du i listrutan Ytfyllning.  
Du kan även förse skrafferingen med en bakgrundsfärg.  
Bitmap  
Ytan fylls med ett bitmap-mönster från den aktuella bitmaptabellen.  
Valet gör Du i listrutan Ytfyllning.  
Du kan definiera ett eget bitmap-mönster eller ladda ett mönster från en pixelgrafikfil och lägga till det på listan.  
Öppna i så fall t ex en %PRODUCTNAME Draw-teckning, rita en rektangel (eller rita rektangeln i ett textdokument med utrullningslisten Ritfunktioner) och öppna sedan dess snabbmeny.  
Välj sedan kommandot Yta...  
Nu kan Du rita eller ladda ett mönster på fliken Bitmapmönster.  
Ytfyllning  
Om Du har valt något av alternativen Färg, Färggradient, Skraffering eller Bitmap, visas motsvarande tabell, där Du kan välja önskad ytfyllning.  
Förutom grundfärger som "magenta" finns även många färgnyanser såsom "blekgul "att välja på.  
Här ser Du även namnet på färgen på ett markerat objekt i en öppet dokument när den färgen inte finns med på den aktuella färgtabellen.  
Om Du vill måla fler objekt med denna nya färg, kan Du i dialogrutan Format - Yta - Färger lägga till den i färgtabellen.  
Steglängd  
Det här området visas bara när Du har valt alternativfältet Färggradient.  
Du kan här välja mellan automatisk och manuell inställning av steglängden.  
automatisk  
Med den här kryssrutan väljer Du automatisk steglängd på färggradienten.  
Steglängd  
Här kan Du ange färggradientens steglängd.  
Följande egenskaper visas bara om alternativfältet Bitmap är valt.  
Storlek  
I det här området definierar du bitmapstorlek.  
Relativ  
Klicka här om du vill förändra bitmapstorleken i förhållande till ytan.  
Om du klickar en gång i rutan, visas måttangivelserna i procent i rotationsfälten Bredd och Höjd.  
Om du klickar en gång till visas angivelserna i måttenheter.  
Original  
Om du vill behålla bitmapmönstrets ursprungliga storlek, markerar du den här rutan.  
Bredd  
Här kan du ändra bitmapmönstrets bredd.  
Höjd  
Här kan du ändra bitmapmönstrets höjd.  
Position  
Här väljer du bitmapmönstrets placering.  
Den aktuella placeringen visas med en röd punkt.  
X-offset  
I det här rotationsfältet kan du förvränga en bitmap i horisontell riktning.  
Y-offset  
I det här rotationsfältet kan du förvränga en bitmap i vertikal riktning.  
Sida vid sida  
Klicka här om Du vill att objektfyllningen ska göras sida vid sida.  
Anpassa  
Med Anpassa anger Du att objektfyllningen ska anpassas till ytans storlek.  
Förskjutning  
I det här området kan du styra förskjutningen av rader eller kolumner i bitmapmönstret.  
Rad  
Välj det här alternativfältet om du vill förskjuta de enskilda raderna i bitmapmönstret.  
Ange förskjutningsmåtten i listrutan intill.  
Kolumn  
Välj det här alternativfältet om du vill förskjuta de enskilda kolumnerna i bitmapmönstret.  
Ange förskjutningsmåtten i listrutan intill.  
Procent  
Här anger Du värdet på rad - eller kolumnförskjutningen i procent.  
Skraffering bakgrund  
Området visas bara när Du har valt Skraffering som typ av ytfyllning.  
Bakgrundsfärg  
För att du ska kunna tilldela en skraffering en bakgrundsfärg måste den här rutan vara markerad.  
Listrutan Bakgrundsfärg  
I den här listrutan väljer du en färg.  
Färger  
Här ställer du in färgen på en yta.  
Det finns mer information om den här fliken i hjälpen till Verktyg - Alternativ - %PRODUCTNAME - Färger.  
Färggradienter  
När du har markerat en yta kan du göra ändringar i en fördefinierad färggradient här eller lägga till nya färggradienter.  
Dessutom kan du ladda eller skapa en ny färggradienttabell.  
Färggradienter som tilldelats ett objekt roterar med när du roterar objektet.  
Typ  
I den här listrutan kan Du välja mellan färggradienttyperna Axialt, Linjär, Radiellt, Ellipsoid, Kvadratisk och Rektangulär.  
Centrum X  
Måttet anges i% av ytans totala bredd.  
Ett värde på 0% innebär att centrum placeras vid vänstra kanten.  
Ett värde på 100% innebär att centrum placeras vid högra kanten.  
Det här alternativet är endast tillgängligt för färggradienttyperna Radiellt, Ellipsoid, Kvadratisk och Rektangulär.  
Centrum Y  
Måttet anges i% av ytans totala höjd.  
Ett värde på 0% innebär att centrum placeras vid den övre kanten.  
Ett värde på 100% innebär att centrum placeras vid den nedre kanten.  
Det här alternativet är endast tillgängligt för färggradienttyperna Radiellt, Ellipsoid, Kvadratisk och Rektangulär.  
Vinkel  
Här anger Du rotationsvinkel för färgradienttyperna Linjär, Axial, Ellipsoid, Kvadratisk och Rektangulär.  
Marginal  
Här anger Du ytandelen för ursprungsfärgen i förhållande till färggradienten.  
Måttet anges i% av totala ytan.  
Ett värde på 100% innebär att färggradienten dämpas ut.  
Från  
Välj en startfärg för färggradienten i listrutan.  
I rotationsfältet kan Du definiera startfärgens intensitet.  
Till  
Välj en slutfärg för färggradienten i listrutan.  
I rotationsfältet kan Du definiera slutfärgens intensitet.  
Färggradienter  
Välj önskad färggradient här.  
Lägg till...  
Med den här kommandoknappen kan Du lägga till en egendefinierad färggradient i den aktuella färggradienttabellen.  
Ange ett namn i dialogrutan Namn.  
Ändra...  
Med den här kommandoknappen ersätter Du inställningarna för en färggradient med de aktuella iinställningarna.  
Välj den färggradient som Du vill ändra i dialogrutan Namn.  
Ladda färggradienttabell  
Med den här ikonen öppnar du dialogrutan Öppna.  
Spara färggradienttabell  
Med den här ikonen öppnar Du dialogrutan Spara som.  
Skrafferingar  
När du har markerat en yta kan du göra ändringar i en fördefinierad skraffering här eller lägga till nya skrafferingar.  
Dessutom kan du ladda eller skapa en ny skrafferingstabell.  
Egenskaper  
I området Egenskaper kan du definiera avstånd och vinkel för skrafferingen.  
Avstånd  
I det här rotationsfältet definierar Du avståndet mellan två skrafferingslinjer.  
Vinkel  
Här definierar Du lutningsvinkeln för skrafferingslinjerna.  
Grafiskt alternativfält  
I det här området kan du välja önskat gradtal direkt.  
Aktuell vinkel är markerad med en röd punkt.  
Linjetyp  
I den här listrutan kan Du välja mellan linjetyperna Enkel, Korsad eller Trippel.  
Linjefärg  
Här väljer Du önskad linjefärg från aktuell färgpalett.  
Tabell  
Du kan skapa egna skrafferingsvarianter med utgångspunkt från de medföljande skrafferingstabellerna.  
Du kan ändra skrafferingar eller lägga till egna skrafferingsutkast.  
Listrutan Skrafferingar  
Här väljer Du önskad skraffering från listan.  
Lägg till...  
Med den här kommandoknappen kan Du lägga till en egendefinierad skraffering i aktuell skrafferingstabell.  
Skapa en ny skraffering genom att ange alternativ på den här fliken och klicka sedan på Lägg till...  
Då visas dialogrutan Namn, där Du kan ange ett namn för den nya skrafferingen.  
Den nya skrafferingen sparas automatiskt.  
Ändra...  
Med den här kommandoknappen kan Du ersätta inställningarna för en skraffering med aktuella inställningar.  
I dialogrutan Namn anger Du namnet för den skraffering som de aktuella inställningarna ska gälla för.  
Ändringen sparas automatiskt.  
Ladda skrafferingstabell  
Med den här ikonen öppnar du dialogrutan Öppna.  
Spara skrafferingstabell  
Med den här ikonen öppnar Du dialogrutan Spara som.  
Bitmapmönster  
När du har markerat en yta kan du här göra ändringar i ett fördefinierat bitmapmönster och lägga till ett nytt pixelmönster.  
Dessutom kan du ladda eller skapa en ny bitmapmönstertabell.  
Mönstereditor  
I detta område med 8x8 pixlar definierar du förgrunds - och bakgrundsfärgen för pixelmönstret och pixelmönstret som sådant.  
Tabell  
Den förinmatade bitmapsmönstertabellen fungerar som utgångspunkt för Dina egna pixelmönstervariationer.  
Du kan ändra pixelmönster och lägga till egna pixelmönsterutkast.  
Förgrundsfärg  
Välj en förgrundsfärg här.  
Bakgrundsfärg  
Välj en bakgrundsfärg här.  
Bitmapsmönster  
Välj önskat bitmapsmönster ur listan i listrutan.  
Lägg till...  
Med denna kommandoknapp kan Du lägga till Dina egendefinierade pixelmönster i den aktuella bitmapsmönstertabellen.  
Namn väljer Du i dialogrutan Namn.  
Ändra...  
Med denna kommandoknapp kan Du skriva över inställningarna för ett pixelmönster med de aktuella inställningarna.  
I dialogrutan Namn väljer Du det pixelmönster som ska ändras.  
Import...  
Dialogrutan Import är identisk med dialogrutan Infoga grafik.  
Ladda bitmaptabell  
Med denna symbol kommer Du till dialogrutan Öppna.  
Spara bitmaptabell  
Med denna ikon öppnar Du dialogrutan Spara som.  
Skugga  
Här bestämmer du om den markerade ytan ska förses med en skugga.  
Med hjälp av Format - (Objekt / Grafik / Tabell) - Inramning definierar Du skuggan för en bild eller ett annat objekt som inte är ett ritobjekt.  
Egenskaper  
Du kan tilldela alla ytor en skugga oberoende av vald ytfyllning.  
Skuggan motsvarar en kopia av den markerade ytan, men är inget självständigt teckningselement.  
Använd skugga  
Aktivera den här rutan om ytan ska ha en skugga.  
Justering  
Här väljer du en position för skuggan.  
Den aktuella positionen visas med en punkt.  
Avstånd  
Ange avståndet mellan skuggan och den markerade ytan eller ställ in avståndet med hjälp av pilknapparna bredvid textfältet.  
Färg  
Här väljer du färg till skuggan.  
Transparens  
Här kan du välja ett transparensvärde för skuggan, mellan 0% (täckande färg) och 100% (osynlig).  
Skugga  
Med den här ikonen på objektlisten aktiverar du respektive inaktiverar skuggan för det markerade objektet.  
Om inget objekt är markerat växlar ikonen till förinställningen Skugga för nya objekt.  
Skugga  
Skugga  
Med den här ikonen aktiverar du respektive inaktiverar du skuggan för det markerade objektet.  
Om inget objekt är markerat, växlar ikonen till förinställningen Skugga för nya objekt.  
Skugga  
Transparens  
Här definierar du om en yta ska visas transparent och med vilken intensitet det ska göras.  
Transparensläge  
I området Transparensläge bestämmer du om och vilken typ av färg som ska visas transparent.  
Ingen transparens  
Om du klickar på det här alternativfältet får den aktiva färgen ingen transparens.  
Den här inställningen är förvald.  
Transparens  
Det här alternativet ger en jämn transparens.  
Rotationsfält Transparens  
I det här rotationsfältet höjer eller sänker du transparensen i det markerade grafikobjektet.  
Fältet är bara aktivt om läget Transparens har aktiverats.  
Värden från 0% (inte allt genomskinlig) till +100% (helt och hållet genomskinlig) är möjliga.  
Gradient  
Om det här alternativet är markerat, kan du välja mellan flera gradienttyper.  
Typerna och deras inställningar hittar du i området Transparensgradient.  
Gradient  
Om det valda transparensläget är en Transparensgradient, kan Du göra mer exakta inställningar i det här området.  
Typ  
I listrutan kan Du välja önskad typ.  
Alternativen är "Lineär", "Radiell", "Axial", "Ellipsoid", "Kvadratisk" och "Rektangulär ".  
Centrum X  
För vissa typer av transparensgradient (t ex Kvadratisk) kan Du här ange med hur många procent centrum för färgförändringen ska förskjutas längs X-axeln.  
Med 100% sker förskjutningen med 50% åt vänster och 50% åt höger.  
Centrum Y  
För vissa typer av transparensgradient (t ex Radiell) kan Du här ange med hur många procent centrum för färgförändringen ska förskjutas längs Y-axeln.  
Med 100% sker förskjutningen med 50% nedåt och 50% uppåt.  
Vinkel  
Du kan ställa in vinkeln på färgförskjutningen genom att ange ett värde mellan 0 ° och 360 ° i den här rotationsrutan.  
Den inställningen kan göras för alla typer.  
Kant  
Om färgförändringen ska vara försedd med en kantlinje, kan Du ange dess storlek i procent här.  
Alltefter den valda typen får Du naturligtvis en särskild kantlinjeeffekt.  
Rotationsfältet kan Du använda för alla typer.  
Startvärde  
Här kan Du ange ett värde på transparensintensiteten i färgförändringens start.  
Det är också det förinställda värdet.  
Slutvärde  
Det kan vara högst 100%.  
Det är också det förinställda värdet.  
Förhandsvisning  
Innan Du bekräftar en inställning eller ändring med OK kan Du se hur den ser ut i den här exempelrutan.  
Text  
Här kan du placera ett text-ritobjekt.  
Rektangeln som omger objektet definierar de kanter som används av funktionerna i denna dialogruta vid justeringen.  
Justera först texten innan Du roterar eller ändrar objektets dimensioner.  
Text  
I detta område anpassar Du texten och ritobjektets ramar till varandra.  
Anpassa bredd till text  
Markera den här rutan om du vill att ramens bredd ska anpassas till textens bredd.  
Anpassa höjd till text  
Markera den här rutan om du vill att ramens höjd ska anpassas till textens höjd.  
Anpassa till ram  
Markera den här rutan om du vill att texten ska anpassas till ramen.  
Textens bredd och höjd skalas så att den exakt fyller ramen.  
Konturflöde  
Markera den här rutan om du vill att konturflödet ska anpassas till texten.  
Avstånd till ram  
I det här området kan du definiera textens avstånd från ritobjektets ram.  
Positiva avstånd krymper texten i motsvarande riktning.  
Du kan också ställa in negativa värden om texten ska fortsätta utanför ramen.  
Vänster  
I detta rotationsfält definierar Du textavståndet från ramens vänsterkant.  
Höger  
I detta rotationsfält definierar Du textavståndet från ramens högerkant.  
Överkant  
I detta rotationsfält definierar Du textavståndet från ramens överkant.  
Underkant  
I detta rotationsfält definierar Du textavståndet från ramens underkant.  
Textförankring  
I det här området definierar du textförankringen.  
Grafiskt alternativfält  
I detta område kan Du definiera den punkt som texten i ramen ska förankras till.  
Denna funktion syns bara när texten inte är dimensionerad att fylla hela ramen.  
Hel bredd  
Om du markerar den här rutan väljer du textförankringen för hela ritobjektets bredd.  
Position och storlek  
Med det här kommandot kan du bl.a. bestämma position och storlek för ett markerat ritobjekt eller kontrollfält.  
Om du har markerat en förklaring heter den här dialogrutan Förklaring.  
Position  
Här definierar du positionen för ett markerat ritelement eller kontrollfält.  
Position  
I det här området definierar du positionen för den markerade objektpunkten.  
Positionen visas med en punkt i det grafiska alternativfältet.  
Om du vill markera en annan objektpunkt klickar du på den önskade positionen.  
Vid roterade eller cirkelformade teckningselement visas stödpunkternas positioner.  
Position X  
Här anger du det vågräta avståndet mellan vänster sidmarginal och den markerade objektpunkten.  
Position Y  
Här anger du det lodräta avståndet från den övre sidmarginalen till den markerade objektpunkten.  
Skydda  
Markera den här rutan om du vill förhindra att objektets ska kunna flyttas från sin aktuella position med musen.  
Baspunkt  
I det här grafiska alternativfältet kan du välja en baspunkt.  
Den valda baspunkten visas med en röd punkt.  
Förankring  
Här bestämmer du var teckningselementet eller kontrollfältet ska förankras.  
Ankare  
I den här listrutan väljer du förankring..  
Position  
Här bestämmer du objektets placering om du har valt förankringen Som tecken.  
Storlek  
Här bestämmer du storleken för ett markerat ritelement eller kontrollfält.  
För 3D-objekt definierar du storleken för aktuell 2D-projektion på papperet.  
Storlek  
I det här området väljer du storleken för det markerade objektet.  
I det grafiska alternativfältet väljer du baspunkten för storleksändringen.  
Den aktuella baspunkten är markerad.  
Baspunktens läge ändras inte när objektets storlek ändras.  
Bredd  
Här anger du bredden för det markerade objektet.  
Höjd  
Här anger du höjden för det markerade objektet.  
Anpassa proportionellt  
Markera den här rutan om storleken på objektet ska förändras proportionellt.  
Skydda  
Markera den här rutan om du vill förhindra att objektets aktuella storlek kan ändras med musen.  
Baspunkt  
I det här grafiska alternativfältet kan du definiera baspunkten.  
Den baspunkt som används för närvarande är markerad med en punkt.  
Anpassa  
I det här området anpassar du objektramens bredd och höjd till motsvarande mått för texten.  
Anpassa bredd till text  
Markera här om du vill att objektramens bredd ska anpassas till textens bredd.  
Anpassa höjd till text  
Markera här om du vill att objektramens höjd ska anpassas till textens höjd.  
Om du klickar här visas det markerade objektet i originalstorlek.  
Rotation  
Här kan du rotera ett markerat ritobjekt genom att välja rotationspunkt och rotationsvinkel.  
Om du väljer en rotationspunkt utanför teckningselementet, kan det hända att teckningselementet inte finns kvar på sidan efter rotationen.  
Rotationspunkt  
Den är markerad med en punkt i det grafiska alternativfältet.  
Du kan flytta den till valfri plats.  
Position X  
Här anger du rotationspunktens vågräta avstånd från den vänstra sidkanten.  
Position Y  
Här anger du rotationspunktens lodräta avstånd från den övre sidkanten.  
Förinställningar  
I det här området kan du välja en av standardrotationspunkterna.  
Den rotationspunkt som för tillfället används visas med en punkt.  
Rotationsvinkel  
I det här området kan du bestämma rotationsvinkeln.  
Vinkel  
Ange rotationsvinkeln i rotationsfältet.  
Förinställningar  
I det här området kan du definiera rotationsvinkeln i steg om 45°.  
Den aktuella vinkeln visas med en punkt.  
Snedställ / hörnradie  
Här kan du snedställa ett ritobjekt som är markerat och i förekommande fall ändra hörnradien.  
Hörnradie  
Det här området är aktivt bara om Du med ritfunktionernas hjälp har skapat ett rätvinkligt hörn.  
Här kan Du runda ett sådant hörn.  
Radie  
I det här rotationsfältet anger Du radien för det markerade hörnet.  
Snedställ  
I det här området kan Du snedställa eller böja ytan.  
Vinkel  
Här anger Du den vinkel med vilken ytan ska böjas.  
Förklaring  
Om du har markerat en förklaring kan du bestämma utseendet för den här.  
Grafiska alternativfält  
Här väljer du typ av förbindelselinje till förklaringen.  
Avstånd  
I det här rotationsfältet anger du avståndet mellan linjen och förklaringen.  
Fäste  
I det här kombinationsfältet väljer du linjens fäste till den markerade förklaringen.  
Beroende på dina val i den här rutan ändras rotationsfältet som finns till höger om den.  
Längd  
I det här rotationsfältet definierar du linjens längd från förklaringen till knicken på en vinklad linje.  
Det här rotationsfältet är bara aktivt om du har valt "Vinklad linje med en knick" och rutan Optimal inte är markerad.  
Optimal  
Klicka här om du vill visa en vinklad linje med en knick optimalt.  
Spegelvänd  
Med det här kommandot kan du spegla ett ritobjekt som är markerat.  
Du kan spegla både horisontellt och vertikalt.  
Det här menykommandot är bara synligt när ett ritobjekt är markerat i ett dokument.  
Vertikalt  
Med det här kommandot spegelvänder du objekt vertikalt.  
Utgångsobjektets överkant blir då det spegelvända objektets underkant.  
Horisontellt  
Med det här kommandot spegelvänder du objekt horisontellt.  
Utgångsobjektets vänstra sida blir då det spegelvända objektets högra sida.  
Placering  
Här sammanfattas de kommandon som används för att lägga objekt "på varandra".  
Den här funktionen kan du bara använda när ett motsvarande objekt är markerat i dokumentet.  
Det kan röra sig om en ram, ett grafikobjekt, ett ritobjekt, ett kontrollfält eller ett annat infogat objekt, t.ex. ett OLE-objekt eller ett diagram.  
Tänk dig att dina sidor består av tre genomskinliga skikt: textskiktet, grafikskiktet i förgrunden och grafikskiktet i bakgrunden.  
Som grafikskikt betecknas här alla skikt som innehåller grafik, teckningar, ramar eller andra objekt.  
De här skikten ligger ovanpå varandra; det ena innehåller texten, de andra grafiken eller andra objekt.  
Alla objekt ligger ovanpå varandra i grafikskiktet med det först ritade grafikelementet eller det först skapade objektet underst och de följande ovanpå, och de överlappar eller täcker då de undre.  
Varje nytt element syns först i förgrundens grafikskikt och täcker alltså textskiktet.  
För kontrollfält till formulär finns dessutom ett kontrollfältsskikt.  
Kontrollfält finns enbart i kontrollfältsskiktet.  
De ritas alltid sist när sidan byggs upp och ligger alltså optiskt sett framför alla andra objekt och texten på sidan.  
Men om du markerar objekt sker det fortfarande efter den interna objektordningen.  
Om du t.ex. först ritar ett kontrollfält och sedan en rektangel, som delvis täcker kontrollfältet, och därefter klickar på det område som kontrollfältet och rektangeln gemensamt upptar på skärmen, så markeras alltid rektangeln.  
Med de första fyra punkterna på undermenyn påverkar du ordningsföljden för grafikelement respektive objekt ovanpå varandra i grafikskiktet, medan de två följande punkterna ordnar in de markerade grafikelementen respektive objekten framför eller bakom textskiktet.  
Längst fram  
Med denna funktion placeras det markerade objektet längst fram.  
Om det redan finns andra objekt på samma ställe täcks det över helt eller delvis.  
Längre fram  
Med detta kommando flyttar du det markerade objektet ett steg längre fram.  
Längre bak  
Med detta kommando flyttar du det markerade objektet ett steg längre bak.  
Längst bak  
Med det här kommandot placerar du det markerade objektet längst bak.  
Om det finns andra objekt på samma ställe kommer det aktuella objektet att döljas helt eller delvis av dessa.  
I förgrunden  
Med detta kommando placerar du ett markerat objekt eller markerade objekt i förgrunden.  
De placeras framför texten och täcker den.  
Den här funktionen är bara tillgänglig om du har markerat ett eller flera ritobjekt.  
Nya ritobjekt visas automatiskt i förgrunden.  
Därför kan du bara använda det här kommandot om du själv har placerat ritobjekten i bakgrunden innan.  
I bakgrunden  
Med kommandot I bakgrunden på snabbmenyn eller med ikonen I bakgrunden placerar du ett markerat ritobjekt i bakgrunden.  
Det placeras och visas bakom texten.  
Ibland kan du inte klicka på och markera ett objekt som du placerat i bakgrunden.  
Då väljer du ikonen Urval på utrullningslisten Ritfunktioner.  
Rita sedan upp en markeringsrektangel runt hela objektet.  
Förankring  
Med förankring kan du välja om det markerade objektet ska förankras vid sidan eller vid cellen vid sidan, vid tecken, som tecken eller vid det markerade stycket.  
Om objektet är inbäddat i en ram kan Du även förankra objektet mot ramen.  
När en ram eller ett bildobjekt skapas, undersöks om objektet finns helt och hållet i en (annan) ram.  
I så fall förankras det till stycket inuti den ramen.  
Vid sidan  
Med detta kommando förankras ett markerat objekt vid sidan.  
Om du ändrar texten kan objektet inte längre flyttas till en annan dokumentsida.  
Ändringar i textområdet påverkar inte ramens placering.  
Om du valt den här förankringen visas ankarsymbolen i det övre vänstra hörnet.  
Vid stycket  
Med det här kommandot förankrar du ett markerat objekt vid aktuellt stycke.  
Om placeringen av det aktuella stycket ändras genom textändringar flyttas även ramen med.  
Om denna förankring är markerad visas ankarsymbolen i högra marginalen i höjd med objektets överkant.  
Vid tecken  
Med det här kommandot förankras ett markerat objekt vid aktuellt tecken.  
Ett objekt som är förankrat vid ett tecken följer med om det tillhörande tecknet flyttas i dokumentet.  
I motsats till förankringen "som tecken" står objektet inte som en bokstav i texten, utan dess horisontala och vertikala placering beräknas med ledning av positionen för det tecken som det är förankrat till.  
Om Du markerar ett objekt som är förankrat till ett tecken, visar en ankarsymbol vilket tecken det gäller.  
För ett objekt som är förankrat till ett tecken kan Du ange placering i förhållande till tecknet.  
Öppna dialogrutan för redigering av objektegenskaper och välj sidan fliken Typ.  
Om Du i området Position anger objektets placering i horisontalled i förhållande till ett tecken, visas ett rött lodrätt streck som referens i förhandsvisningsfältet.  
Det strecket motsvarar det blinkande markörstrecket när detta befinner sig framför det tecken som Du har angett som ankare.  
Vid cellen  
Med det här kommandot kopplas teckningselementets ankarpunkt till cellen.  
Teckningselementet är knutet till cellen.  
Om du väljer den här förankringen, visas ankarsymbolen i höjd med teckningselementets övre vänstra hörn.  
Vid ram  
Med detta kommando förankras ett markerat objekt vid ramen som omger objektet.  
Den här funktionen är bara tillgänglig för objekt som är infogade i en ram.  
Som tecken  
Med detta kommando förankrar du ett markerat objekt som tecken.  
Ett objekt som förankrats som tecken står som en normal bokstav i texten och påverkar därför radhöjd och brytning.  
Då texten ändras i stycket flyttas också objektet i sidled.  
Redigera punkter  
Med den här funktionen kan du redigera punkterna i ett markerat ritobjekt.  
Med ikonen Redigera punkter på Objekt - eller Alternativlisten Objekt - eller Alternativlisten Objektlisten sätter du på eller stänger av redigeringsläget.  
Du kan också välja kommandot Redigera punkter via snabbmenyn till ett markerat ritobjekt.  
Du kan också välja kommandot Redigera punkter via snabbmenyn till ett markerat ritobjekt.  
Om redigeringsläget är aktiverat, kan du flytta varje punkt på en kurva med musen.  
Dessutom kan du flytta punkterna som används för att definiera en polygon.  
Det finns fler ikoner för hantering av punkter på Bézierobjektlistan.  
FontWork  
FontWork används för utformning av teckeneffekter.  
De här effekterna kan du tilldela textobjekt som du har skapat med hjälp av ritfunktionerna på verktygslisten (ikonen Visa ritfunktioner).  
Med FontWork kan du justera ett markerat textobjekt till "osynliga" halvcirklar, cirkelbågar, cirklar och till frihandslinjer.  
Du kan när som helst ersätta justeringsobjektet med ett annat justeringsobjekt.  
Menykommandot FontWork hittar du på menyn Format när du har markerat ett textritobjekt i ett dokument.  
Funktionerna i FontWork-fönstret kan bara användas för textobjekt.  
Justeringsikoner  
I det här området kan du tilldela en markerad text formen av en halvcirkel, cirkelbåge eller sluten cirkel genom att välja en av de många ikonerna.  
I den övre delen av FontWork finns det olika symboler.  
Om du klickar på någon av dem kommer den markerade texten i dokumentet att justeras på motsvarande sätt.  
I den övre raden finns ikoner för olika halvcirklar.  
Här väljer du bland justeringstyperna Övre halvcirkel, Undre halvcirkel, Vänster halvcirkel och Höger halvcirkel.  
Halvcirklar  
Därefter finns ikoner för olika cirkelbågar.  
Här väljer Du mellan de olika justeringsalternativen Övre cirkelbåge, Undre cirkelbåge, Vänster cirkelbåge och Höger cirkelbåge.  
Cirkelbågar  
Till sist kan Du också välja mellan olika cirkeljusteringsalternativ:  
Öppen cirkel, Stängd cirkel, Stängd cirkel II och Öppen cirkel lodrätt.  
Cirklar  
Om Du klickar på ikonen Av tar Du bort anpassningen av textobjektet till justeringsobjektet.  
Av  
Med symbolen Rotera roterar Du textobjektets tecken så att de står med sin bas på justeringsobjektets konturlinje.  
Rotera  
Textobjektet följer justeringsobjektets konturlinje.  
Upprätt  
Med ikonen Tippa horisontellt tippas textobjektets tecken horisontellt.  
Tippa horisontellt  
Med ikonen Tippa vertikalt tippas textobjektets tecken vertikalt.  
Tippa vertikalt  
Om Du klickar på Löpriktning vänds textens aktuella löpriktning.  
Textobjektet placeras då inte ovanför utan under justeringsobjektets konturlinje.  
Löpriktning  
Om du klickar på Vänsterjusterat placeras textobjektet till vänster i justeringsobjektet.  
Vänsterjusterat  
Om du klickar på Centrerat placeras textobjektet i mitten av justeringsobjektet.  
Centrerat  
Om du klickar på Högerjusterat placeras textobjektet till höger i justeringsobjektet.  
Högerjusterat  
Med ikonen AutoTextstorlek ändrar du textobjektets teckenstorlek så att textobjektet upptar hela konturlinjen.  
AutoTextstorlek  
Ange i rotationsfältet Avstånd avståndet mellan justeringselementet och baslinjen för de enskilda tecknen.  
Avstånd justeringselement - baslinje tecken  
Ange i rotationsfältet Indrag avståndet mellan början på justeringsobjektets konturlinje och textens början.  
Avstånd konturlinje - textbörjan  
Med ikonen Kontur slår Du på och stänger av konturlinjen för det aktuella justeringsobjektet.  
Kontur  
Med ikonen Bokstavskontur slår Du på och stänger av konturlinjen för enskilda tecken i textobjektet.  
Bokstavskontur  
Klicka på skuggikonen Av om tecknen ska visas utan skugga.  
Ingen skugga  
Klickar Du på ikonen Lodrätt kommer tecknen att förses med en lodrät skugga.  
Avståndet mellan tecknet och skuggan anger Du i de båda undre rotationsfälten.  
Lodrätt  
Klickar Du på ikonen Tippa kommer tecknen att förses med en tippad skugga.  
Tippvinkeln och skuggstorleken, som hänför sig till originalstorleken på tecknet, anger Du i de båda undre rotationsfälten.  
Tippa  
Horisontellt avstånd  
I rotationsfältet Avstånd X definierar Du det horisontella avståndet mellan skuggan och tecknet.  
Avstånd X  
Vertikalt avstånd  
I rotationsfältet Avstånd X definierar Du det vertikala avståndet mellan skuggan och tecknet.  
Avstånd Y  
Skuggans färg  
I denna listruta väljer Du en färg på skuggan från den aktuella färgtabellen.  
Grupp  
I den här undermenyn hittar du alla funktioner för gruppering av objekt.  
Arbeta med grupper  
Gå in i grupp:  
Via kommandon i menyn eller snabbmenyn, via F3 eller genom att dubbelklicka på en grupp.  
I gruppen är först inget objekt markerat.  
Inom en grupp:  
Alla objekt, som inte hör till gruppen som du har gått in i, visas med svagare färger (ghosted).  
Navigering mellan objekten i en grupp: med hjälp av Tab och Skift+Tab växlar du fram och tillbaka mellan objekten.  
Lämna grupp: via menykommando eller Ctrl+F3 eller genom att dubbelklicka bredvid alla objekt.  
När du lämnat gruppen är den markerad.  
Gruppera  
Upphäv gruppering  
Gå in  
Lämna  
Gruppering / Gruppera  
Med det här kommandot sammanför du markerade objekt till en grupp.  
Därvid behåller de enskilda elementen sina egna egenskaper.  
Genom att skapa grupper kan Du förhindra att de inbördes förhållandena mellan elementen i fråga ändras.  
Du kan dessutom sammanföra flera grupper till en ny (överordnad) grupp.  
Upphäv gruppering  
Med det här kommandot upphäver du den markerade grupperingen.  
Upphäv gruppering påverkar bara en nivå hos de sammanfattade elementen.  
Om gruppen innehåller fler undergrupper där du vill upphäva grupperingen, måste du göra det i ett separat arbetssteg.  
Gå in i gruppering  
Med detta kommando kommer du till den första nivån i grupphierarkin för det markerade gruppobjektet.  
Där kan du markera och redigera de sammanfogade elementen var för sig.  
Gruppobjektets gruppering upphävs inte genom denna åtgärd.  
Du kan gå in i en gruppering genom att dubbelklicka på ett objekt i gruppen.  
Som optiskt svar visas sedan blekare färger på alla andra objekt och grupper som inte hör till den grupp som du gick in i.  
Senare kan du lämna gruppen genom att dubbelklicka utanför gruppens begränsningsrektangel.  
När du har lämnat gruppen förblir den markerad i sin helhet.  
Om du klickar på ett gruppobjekt och samtidigt håller ner Kommando Ctrl -tangenten, så markeras bara det delobjekt som du klickade på, utan att du behöver välja kommandot Gå in i gruppering.  
Detta är bekväma möjligheter att redigera grupperingar utan att behöva använda kommandot Gå in i gruppering.  
Lämna gruppering  
Med det här kommandot kan Du avsluta redigering av de enskilda objekten i ett gruppobjekt.  
För gruppobjekt som innehåller underliggande gruppobjekt kommer Du till närmast högre nivå med det här kommandot.  
Löptext  
Här förser du ett textritobjekt med effekter.  
Effekter animerad text  
I det här området finns alla element som du behöver för att skapa en texteffekt.  
Effekt  
I den här listrutan finns alla effekter som kan väljas:  
Ingen effekt, Blinka, Genomlöpa, Löpa fram och tillbaka, Löpa in i.  
Du kan inte använda symbolknapparna om du väljer Ingen effekt eller Blinka.  
Åt vänster  
Om du klickar på den här symbolen kommer texten som står i ritobjektet att löpa från höger till vänster.  
Åt vänster  
Åt höger  
Om du klickar på den här symbolen kommer texten som står i ritobjektet att löpa från vänster till höger.  
Åt höger  
Uppåt  
Om du klickar på den här symbolen kommer texten att löpa nedifrån och upp.  
Uppåt  
Nedåt  
Om du klickar på den här symbolen kommer texten att löpa uppifrån och ned.  
Nedåt  
Egenskaper  
Text synlig vid start  
Om du markerar det här fältet syns texten redan när du startar effekten.  
Om du har valt effekten Löpa in i kan du inte välja det här alternativet.  
Text synlig vid avslutning  
Om du markerar det här fältet syns texten när du avslutar effekten.  
Om du har valt effekten Löpa in i kan du inte välja det här alternativet.  
Antal  
I det här området definierar du antalet upprepningar.  
Kontinuerligt  
Om den här rutan är markerad upprepas den valda effekten hela tiden.  
Om du bara vill upprepa effekten några gånger avmarkerar du Kontinuerligt och anger det önskade antalet repetitioner i rotationsfältet.  
Kontinuerligt  
I det här rotationsfältet definierar du antalet gånger som effekten ska upprepas.  
Steglängd  
I det här området definierar du effektens steglängd.  
Pixel  
Om Pixel har markerats (standardinställning) är steglängden definierad i måttenheten pixel.  
Om du avmarkerar Pixel anges steglängden i centimeter i rotationsfältet.  
Pixel  
I rotationsfältet ändrar du pixelantalet.  
Fördröjning  
I det här området definierar du effektens hastighet.  
Automatisk  
Om Automatisk är markerad upprepas effekten med en hastighet som är definierad av programmet.  
Om du själv vill bestämma hastigheten avmarkerar du Automatisk och anger fördröjningen i rotationsfältet.  
Automatisk  
Ju större värde du anger desto längre blir fördröjningen.  
Radhöjd  
Här kan du ändra de markerade radernas radhöjd.  
Du kan även ställa in radhöjden genom att dra mellanrummet mellan radrubrikerna; i detta fall visas den aktuella radhöjden i tipshjälpen.  
Om Du dubbelklickar på mellanrummet ställer Du in den optimala radhöjden för raden ovanför mellanrummet.  
Höjd  
I detta rotationsfält anger Du den önskade radhöjden.  
Standardvärde Automatiskt  
Om du markerar den här rutan anpassas radhöjden automatiskt till det använda teckensnittet.  
Om den här rutan är markerad, spärras rotationsfältet Höjd.  
Kolumnbredd  
Här ställer du in bredden för de markerade kolumnerna.  
Då visas bredden i en tipshjälpruta.  
Om Du dubbelklickar på mellanrummet ställs optimal kolumnbredd in för spalterna till vänster om mellanrummet.  
Du kan även ställa in kolumnbredden genom att dra i kolumnlinjerna mellan kolumnhuvudena.  
Genom att dubbelklicka på ett spalthuvud ställer Du in optimal bredd för den tillhörande kolumnen, vilket innebär att den anpassas till kolumninnehållet.  
Bredd  
I det här rotationsfältet kan du ändra bredden på en eller flera kolumner som är markerade i tabellen.  
Standardvärde Automatiskt  
Här ställer Du in kolumnbredden efter bredden på kolumnrubriken.  
Justering  
Dessutom definierar du avståndet till gitterlinjerna, textflödet och skrivriktningen här.  
Du kan alltså placera cellinnehållet i cellen efter dina önskemål.  
Du kan ändra cellinnehållet i horisontell och vertikal riktning och ställa in avståndet till gitterlinjerna.  
Horisontell  
I det här kombinationsfältet kan du ställa in justeringen av cellinnehållet i horisontell riktning.  
Standard  
Med det här alternativet kan du välja den horisontella standardinställningen för cellinnehåll.  
Om Du har markerat alternativet Standard blir siffrorna högerjusterade och texten vänsterjusterad.  
Vänster  
Med det här alternativet vänsterjusterar du innehållet i den markerade cellen.  
Höger  
Med det här alternativet högerjusterar du innehållet i den markerade cellen.  
Centrerat  
Med det här alternativet centrerar du cellinnehållet horisontellt.  
Marginaljustering  
Med det här alternativet marginaljusterar du cellinnehållet.  
Indrag  
Välj hur stort indraget ska vara.  
Med ikonerna Minska indrag och Öka indrag på objektlisten kan du flytta cellinnehållet med det avstånd som du har angett här.  
Vertikalt  
Här kan du justera cellinnehåll vertikalt.  
Standard  
I det här alternativfältet kan Du välja standardinställningen för den vertikala justeringen av cellinnehållet.  
Uppe  
Här justeras cellinnehållet vid cellens övre kant.  
Nere  
Här justeras cellinnehållet mot cellens nedre kant.  
Mitten  
Med det här alternativet centreras cellinnehållet vertikalt.  
Skrivriktning  
I det här området definierar du skrivriktningen för cellinnehållet.  
Med hjälp av den runda kommandoknappen ställer du in skrivriktningen steglöst med musen.  
Om du klickar på den rektangulära kommandoknappen, visas cellinnehållet i vertikal skrivriktning.  
Vinkel  
I rotationsfältet anger du rotationsvinkeln.  
Referenskant  
Med hjälp av de här rutorna definierar du cellinnehållets referenskant.  
Den aktuella positionen för den roterade texten bestäms dessutom av områdena Horisontell och Vertikal.  
Textutsträckning från undre cellkanten.  
Den roterade texten skrivs från den undre kanten.  
Textutsträckning från övre cellkanten.  
Den roterade texten skrivs från den övre kanten.  
Textutsträckning bara inuti cellen.  
Den roterade texten skrivs bara inuti cellen.  
Avstånd till gitterlinjer  
Välj avståndet till gitterlinjerna med rotationsfälten.  
Vänster  
I det här rotationsfältet kan Du ställa in cellinnehållets avstånd till vänster gitterlinje.  
Höger  
I det här rotationsfältet kan Du ställa in cellinnehållets avstånd till höger gitterlinje.  
Överst  
I det här rotationsfältet kan Du ställa in cellinnehållets avstånd till den övre gitterlinjen.  
Underst  
I det här rotationsfältet kan Du ställa in cellinnehållets avstånd till den nedre gitterlinjen.  
Textflöde  
Här definierar Du textflödet i cellen.  
Radbrytning  
Om du markerar den här rutan tillåts automatisk radbrytning i cellkanten.  
Oberoende av det kan du alltid göra en manuell radbrytning med Kommando Ctrl +Retur.  
Avstavning aktiv  
Här aktiverar du avstavningen.  
Avstavningen fungerar i celler och ritobjekt om du har aktiverat radbrytning eller textjustering - horisontell - marginaljustering under den här fliken.  
Arbeta med databastabeller  
Här hittar du hjälp till hur du använder databastabeller.  
Om en tabell har öppnats i utkastläge kan den inte öppnas i datakällvyn.  
Stäng först utkastvyn eller inaktivera redigeringsläget där.  
Datakällvyn  
I datakällvyn är redigeringskommandon tillgängliga på databaslisten och på snabbmenyerna.  
I nedre kanten av datavyn finns en Navigationslist som du använder för att snabbt kunna navigera inom dataposterna.  
Markering i datakällvyn  
I datakällvyn ser du dataposterna i den laddade databastabellen.  
Du kan flytta den här pekaren med piltangenterna uppåt och nedåt eller med kommandoknapparna i fönstrets nedre kant eller genom att klicka med musen på en annan datapost.  
I datakällvyn kan du redigera fält, dataposter eller kolumner på olika sätt.  
Du måste först tala om för %PRODUCTNAME Base vad du vill redigera genom att markera elementen.  
Följande tabell ger en överblick över hur du kan markera olika element i datakällvyn:  
Uppgift  
Åtgärd  
Markera en datapost  
Klicka på radhuvudet  
Markera flera dataposter eller upphäva markering  
Håll ner Ctrl - eller skifttangenten och klicka på radhuvudena  
Markera en kolumn  
Klicka på kolumnhuvudet  
Markera ett enstaka datafält  
Klicka i datafältet  
Markera hela tabellen  
Klicka i det vänstra, övre hörnet  
Redigera tabeller  
Om du ska redigera tabellen (lägga till, ändra eller radera data) kan du använda ikonerna på funktionslisten (Redigera, Spara och Ångra).  
När en %PRODUCTNAME databastabell öppnas skrivskyddad, klickar du först på ikonen Redigera fil på funktionslisten eller på databaslisten, så att tabellen friges för redigering.  
I redigeringsläget kan du t.ex. lägga till nya dataposter och ändra eller radera befintliga data.  
Du kan inte ändra databastabellens struktur, t.ex. datafältens ordningsföljd eller egenskaper, i datavyn.  
Det gör du i tabellutkastet.  
När Du redigerar en sökning övertas ändringarna omedelbart av den tillhörande databastabellen.  
Du kan bara lägga till, ändra eller radera data när sökningen enbart avser en tabell.  
En sökning i flera tabeller öppnas alltid skrivskyddad och kan bara redigeras i sökningsutkast.  
Databastabeller, som behöver ett entydigt index eller en primärnyckel för att entydigt kunna identifiera dataposterna, kan inte redigeras när det inte finns varken index eller primärnyckel i tabelldefinitionen.  
I det här fallet kan du inte skriva in, ändra eller radera data.  
Klippa ut, kopiera, klistra in data  
När du har markerat ett enskilt datafält blir funktionerna Klipp ut, Kopiera och Klistra in tillgängliga.  
Du kan klippa ut eller kopiera innehållet i en tabellcell för att sedan infoga innehållet från urklippet igen i en annan tabellcell.  
Du kan också använda tangentkombinationerna Kommando Ctrl +X, Kommando Ctrl +C respektive kommando Ctrl +V.  
Kopiera med dra-och-släpp i tabellen  
Du kan kopiera fältinnehållet i en tabell med dra-och-släpp.  
Då markerar du helt enkelt innehållet i ett datafält och drar det med musen till ett annat datafält.  
Kopiera mellan tabell och dokument med dra-och-släpp  
Du kan dra vanlig text från ett valfritt %PRODUCTNAME -dokument och släppa den i enskilda celler i en tabell.  
Om det redan finns text i datafältet skrivs den över.  
Markera först datafältet, som texten ska överföras till, i databastabellen.  
Markera sedan den text som ska kopieras i det andra dokumentet och dra den med musen till datafältet som du markerade i steg 1.  
Om tabellen eller sökningen visas i datakällvyn drar du helt enkelt texten från det aktuella dokumentet till datakällvyn.  
En förutsättning för att det ska gå att kopiera texten med dra-och-släpp till en tabell är att tabellen redan är i redigeringsläge.  
Dessutom måste du först markera cellen som texten ska kopieras till.  
Att kopiera genom att dra och släppa från ett %PRODUCTNAME -dokument är bara möjligt med "vanlig" text, vilket innebär att bara alfanumeriska tecken (tecken eller tal) är tillåtna.  
Ja / nej-fält, binär-, bild - och räknare-fält.  
I omvänd riktning kan du också kopiera data från en databastabell till ett dokument med dra-och-släpp.  
Metoden beskrivs i hjälpen till datakällvyn.  
Navigation inom tabellen  
Om du vill hoppa till olika dataposter kan du använda navigationslisten under datavyn.  
Första dataposten  
Med denna kommandoknapp sätter Du pekaren på den första dataposten.  
Förra dataposten  
Med denna kommandoknapp sätter Du pekaren på förra dataposten.  
Datapostnummer  
Här ser Du numret på den datapost som pekaren i vänster fönsterkant pekar på.  
Här kan Du skriva in ett nummer och trycka på retur, så flyttar Du pekaren direkt till den nya positionen.  
Här visas det totala antalet dataposter som har laddats.  
En stjärna (*) visar att inte alla dataposter har laddats.  
Nästa datapost  
Med denna kommandoknapp sätter Du pekaren på nästa datapost.  
Sista dataposten  
Med denna kommandoknapp sätter Du pekaren på den sista dataposten.  
Ny datapost  
Om du klickar på stjärnsymbolen hoppar insättningspunkten till slutet av databastabellen och du kan mata in en ny datapost här.  
Den här funktionen är bara tillgänglig när databasen är i redigeringsläge.  
Ikonen Redigera på databaslisten eller funktionslisten måste vara intryckt.  
Markering / totalt  
Här visas i formen x / y hur många dataposter som är markerade (x) och hur många det finns totalt (y).  
Om dataposterna håller på att läsas in och räknas i bakgrunden visas i stället för det totala antalet dataposter ett frågetecken (y =?).  
Utformning av tabeller  
På rad - och kolumnhuvudenas snabbmenyer hittar du olika kommandon, med vars hjälp du kan ändra tabellens utseende.  
Du behöver inte spara dina ändringar eftersom %PRODUCTNAME automatiskt övertar ändringarna.  
Om du stänger tabellen och öppnar den igen kan du se att samtliga attribut som du har angett fortfarande gäller.  
Det finns följande kommandon för tabellutformning:  
Tabellformatering  
Radhöjd...  
Kolumnformatering...  
Kolumnbredd...  
Tabellformatering  
Här kan du göra formateringar som gäller för de valda raderna.  
Radera rader  
Med det här kommandot raderar du den aktuella raden eller alla markerade rader efter en kontrollfråga.  
Det här kommandot kan du bara använda om du har klickat på ikonen Redigera på databaslisten eller funktionslisten.  
Fältformatering  
Här kan du formatera den aktuella kolumnen eller de markerade kolumnerna.  
Om du ändrar fältformateringar här påverkar det inte de verkliga formaten för enstaka fält i databasen.  
Här kan Du t ex inte konvertera ett textfält till ett numeriskt fält eller tvärtom.  
De formateringar Du gör här är endast till för visningen.  
Format  
Dölj fält  
Med det här kommandot döljer du det markerade fältet.  
Visa alla fält  
Med det här kommandot visar du alla fält igen som du tidigare har dolt med kommandot Dölj fält.  
Du kan bara välja det här kommandot om alla fält verkligen är dolda.  
3D-effekter  
Här kan du definiera diverse effekter för tredimensionella objekt.  
Du når de olika områdena i det här fönstret via symbolerna i fönstrets övre del.  
Du kan kombinera valfria 3D-objekt till grupper (scener), men ändå kan alla objekt var för sig redigeras, flyttas, kopieras, raderas och så vidare.  
Markera med musen de objekt som ska grupperas och välj sedan Gruppera i snabbmenyn.  
Därefter har du tillgång till kommandona Lämna gruppering, Gå in i gruppering och Upphäv gruppering.  
Du kan även utföra de här åtgärderna via kortkommandon.  
Du kan även utföra de här åtgärderna via kortkommandon.  
Favoriter  
Här kan du se och välja favoriterna.  
Du öppnar det här området via symbolen Favoriter.  
Favoriter är kombinerade egenskaper för 3D-objekt vilka du kan tilldela andra 3D-objekt genom att klicka med musen.  
Favoriter  
Bilderna i favoriterna är identiska med de grafiska objekten som du hittar i Gallery -temat 3D.  
Om du utökar Gallery-temat 3D med ytterligare grafiska objekt, så visas de också under "Favoriter".  
Favoriter  
I det här området väljer du en favorit.  
Markera först ett 3D-objekt i dokumentet och dubbelklicka sedan på favoriterna.  
De är indelade i grupper:  
De ändrar bara det markerade objektets belysning.  
Den första ringen återställer standardbelysningen, utan att göra några andra ändringar.  
Sedan följer några klot som ändrar det markerade objektets textur.  
De fyra stora bokstäver står för extrusionsobjekt.  
Med dem tilldelas det markerade objektet olika 3D-effekter.  
Tilldela bara 3D-attribut  
Med denna kommandoknapp tilldelar du det markerade objektet bara attributen för 3D.  
Tilldela bara 3D-attribut  
Tilldela alla attribut  
Om du vill tilldela det markerade objektet alla attribut väljer du den här kommandoknappen.  
Tilldela alla attribut  
Uppdatera  
Om du klickar här, visar dialogrutan alla egenskaper för det markerade objektet.  
Uppdatera  
Tilldela  
Klicka här om du vill tilldela det markerade objektet de egenskaper som visas i dialogrutan.  
Tilldela  
Omvandla till 3D  
Med den här ikonen omvandlar du ett markerat 2D - till ett 3D-objekt.  
Men en grupp av 2D-objekt kan inte omvandlas till 3D - upphäv först grupperingen.  
Omvandla till 3D  
Omvandla till rotationsobjekt  
Med den här kommandoknappen omvandlar du ett markerat 2D-objekt till ett 3D-rotationsobjekt.  
Men en grupp av 2D-objekt kan inte omvandlas till 3D - upphäv först grupperingen.  
Omvandla till rotationsobjekt  
Perspektiv på / av  
Klicka på denna kommandoknapp för att sätta på eller stänga av den perspektiviska visningen.  
Perspektiv på / av  
Geometri  
Här kan du göra olika inställningar som ändrar ditt objekts geometriska struktur.  
Geometri  
Geometri  
I det här området kan du ändra ett objekts geometri.  
Ett extrusionsobjekt bildas om en framsida dras till den tredje dimensionen på en bana som står lodrätt till framsidan och vars längd anges med värdet Djup.  
Om värdet för djupskalningen inte är lika med 100%, så blir baksidan större eller mindre än framsidan.  
Ett rotationsobjekt uppstår om en 2D-yta roteras runt en axel som ligger på ytans nivå.  
Ytan roteras på en cirkelformig bana till den tredje dimensionen.  
Ett rotationsobjekt har inget värde för Djup, men det kan ha ett värde för Djupskalning.  
Om värdet för slutvinkeln är exakt 360 grader, så ligger framsidan direkt på rotationsobjektets baksida.  
Rundade kanter  
I detta rotationsfält bestämmer Du hur mycket ett objekts kanter ska rundas.  
De 3D-objekt som medföljer programmet, som t ex kuben, kan inte ändras.  
Dra upp en 2D-rektangel och omvandla den med kommandoknappen Omvandla till 3D till en parallellepiped.  
Nu kan Du ändra kanternas rundning.  
Djupskalning  
Detta värde definierar skalningen mellan fram - och baksida hos ett 3D-objekt.  
Baksidan förstoras eller förminskas i förhållande till framsidan med den nämnda procentsatsen.  
Om du t.ex. använder en djupskalning på 10% på en 3D-cylinder, så ser du nu en hård övergång på det ställe där baksidan och framsidan möts.  
Du ser dessutom på vilket sätt cylindern har konstruerats.  
Detta blir ännu tydligare om du i det följande rotationsfältet förminskar slutvinkeln till t.ex. 270 grader.  
Slutvinkel  
I detta rotationsfält ställer Du in vinkeln om 3D-objektet har skapats genom rotation.  
Ifall Du här t ex för en ring anger mindre än 360 grader så visas den som ett mer eller mindre öppet objekt.  
Djup  
I detta rotationsfält bestämmer Du objektets tredimensionella djup i cm.  
Inställningen träder i funktion om Du t ex med kommandoknappen Omvandla till 3D har omvandlat ett 2D-objekt till ett 3D-objekt.  
Segment  
Här anger Du hur många segment som ska användas för att bygga upp ett 3D-objekt.  
Tack vare denna inställningsmöjlighet är det t ex mycket enkelt att omvandla en torus till en tredimensionell triangel genom att Du ställer in antalet 3 för de horisontella segmenten.  
Horisontell  
I detta rotationsfält anger Du antalet vågräta segment.  
Vertikal  
I detta rotationsfält anger Du antalet lodräta segment.  
Normaler  
I det här området finns det fler kommandoknappar som används till att förändra det markerade objektets geometri.  
Objektspecifik  
Med detta alternativ visas objektet på ett anpassat sätt, t.ex. visas ett sfäriskt objekt och rundade områden på ett objekt genom en sfärisk projektion, ett rätvinkligt objekt och platta områden genom en platt projektion.  
Objektspecifik  
Platt  
Välj denna kommandoknapp om rundade former ska visas som små ytor (polygoner).  
Ifall Du samtidigt vill använda läget Flat (platt) på fliken Visning, bör Du ta hänsyn till att i detta fall geometrin Platt används på det aktuella objektet.  
Platt  
Sfärisk  
Med detta alternativ tvingar Du fram en sfärisk visning.  
Sfärisk  
Omvända normaler  
Med detta alternativ omvänds belysningsförhållandena för objektet, så att objektet till synes belyses "inifrån" i stället för utifrån.  
Denna effekt syns bara i öppna 3D-objekt.  
Omvända normaler  
2-sidig belysning  
Hos öppna 3D-objekt definierar Du här en likadan inre och yttre belysning.  
Ifall Du samtidigt har aktiverat Omvända normaler, så belyses objektet bara av omgivningsljuset.  
2-sidig belysning  
Dubbelsidig  
Ifall denna kommandoknapp är aktiverad, så visas 3D-objektet över sitt totala omfång som slutet objekt.  
Denna funktion verkar på 3D-objekt som t ex har skapats genom extrusion ur en fylld frihandslinje som korsar sig själv.  
På grund av 2D-linjens korsning uppkommer vid extrusionen till 3D flera delobjekt.  
Ifall funktionen Dubbelsidig har tilldelats, så har alla delobjekt till 3D-objektet fullständiga botten-, topp - och sidytor.  
Ifall denna funktion inte har aktiverats, så är bara det första delobjektet fullständigt stängt, de andra delobjekten är delvis öppna.  
Dubbelsidig  
Visning  
Här ställer du in hur objekt ska visas.  
Visning  
Visning  
I det här området bestämmer du hur objektet ska visas.  
Läge  
Med de tre lägena Flat, Phong och Gouraud bestämmer du bildskärmsvisningens kvalitet genom att välja en beräkningsmetod.  
Från Flat via Phong till Gouraud ökar visningens kvalitet, men även laddningstiden blir längre.  
Skugga  
Med denna kommandoknapp aktiverar eller inaktiverar Du 3D-skuggan.  
3D-skugga på / av  
Papperslutning  
I detta rotationsfält kan Du ställa in lutningen på den tänkta pappersytan på vilken objekt-skuggan faller.  
Välj bland vinklar från 0 till 90 grader.  
Kamera  
I detta område gör Du inställningar som motsvarar inställningarna för en kamera.  
Avstånd  
I detta rotationsfält kan Du ändra avståndet mellan betraktaren och mitten på ett objekt.  
Brännvidd  
Här ställer Du in med vilken brännvidd objektet ska betraktas.  
Ju mindre brännvidden är desto större blir "fisköge-effekten" som uppstår, medan stora brännvidder motsvarar en "tele-effekt ".  
Belysning  
Här kan du välja och ställa in ljuskällor.  
Du öppnar det här området via symbolen Belysning.  
Belysning  
Belysning  
I detta område väljer Du ljuskällorna och ställer in RGB-värdena samt omgivningsljuset.  
Du kan välja bland åtta ljuskällor som kan definieras fritt.  
Ljuskälla  
Klickar Du en gång till på ikonen så sätts ljuskällan på, klickar Du på nytt så stängs den av.  
När du har markerat ett nytt objekt genom att klicka på det med musen, används den andra ljuskällan om du inte ändrar det.  
Den andra ljuskällan skapar i motsats till den första ljuskällan inte någon högdager och därför förfalskas färgerna inte.  
Ljuset är på  
Ljuset är släckt  
Färgurvalsfält  
I detta urvalsfält väljer Du den aktuella ljuskällans färg.  
Färgernas intensitet har redan tagits hänsyn till.  
Välj färg via färgdialogen  
Omgivningsljus  
Här bestämmer du färgen på omgivningsljuset.  
Omgivningsljuset kan du t.ex. använda när objekt som är för mörka ska göras ljusare.  
Färgurvalsfält  
I detta urvalsfält väljer Du omgivningsljusets färg.  
Välj färg via färgdialogen  
Förhandsvisning  
Det här fönstret används förutom till förhandsvisning av ändringar även för placering av de olika belysningskällorna.  
Du kan med musen justera ljuskällor på en sorts lampram.  
För finjustering använder du fönstrets bildrullningslister.  
Du kan tilldela var och en av ljuskällorna en annan färg.  
Texturer  
Här kan du ändra återgivningen av texturer.  
Du tilldelar ett objekt en textur genom att t.ex. dra en bitmap från Gallery till objektet samtidigt som du håller ner Skift+Ctrl.  
Texturer  
Texturer  
I detta område väljer Du olika inställningar för texturer.  
Typ  
Här kan Du välja mellan visning i svartvit och i färg.  
Svartvit  
Med denna kommandoknapp kan Du tilldela svartvit till texturer.  
Svartvit  
Färg  
Denna kommandoknapp ger en textur i färg.  
Färg  
Läge  
Här bestämmer Du om bara textur ska tilldelas eller textur med andra effekter.  
Bara textur  
Här väljer Du att bara textur ska användas.  
Bara textur  
Textur och skugga  
Här väljer Du att textur och skugga ska användas.  
Textur och skugga  
Projektion X  
Med de tillhörande kommandoknapparna bestämmer Du för Ditt objekts X-axel hur texturen ska placeras.  
Objektspecifik  
Detta alternativ ger en textur som anpassas optimalt till objektet.  
Objektspecifik  
Parallell  
Med detta alternativ skjuts texturen på sätt och vis genom objektet.  
Parallell  
Cirkelformad  
Med denna kommandoknapp läggs texturen sfäriskt runt objektet.  
Cirkelformad  
Projektion Y  
Med de tillhörande kommandoknapparna bestämmer Du för Ditt objekts Y-axel hur texturen ska placeras.  
Objektspecifik  
Detta alternativ ger en textur som anpassas optimalt till objektet.  
Objektspecifik  
Parallell  
Med detta alternativ skjuts texturen på sätt och vis genom objektet.  
Parallell  
Cirkelformad  
Med denna kommandoknapp läggs texturen sfäriskt runt objektet.  
Cirkelformad  
Filtrera  
Med detta alternativ kan Du förbättra objektets utseende.  
Filtrera på / av  
Med denna kommandoknapp kan Du sätta på eller stänga av filterfunktionen.  
Filtrera på / av  
Material  
Här kan du tilldela objekt färger som ser ut som vissa material.  
Du öppnar det här området via symbolen Material.  
Material  
Material  
I detta område kan Du välja olika inställningar som ger Ditt objekt ett visst utseende (t ex träliknande eller metalliskt).  
Favoriter  
Här kan du välja en yta.  
Objektfärg  
I den här listrutan väljer du objektets färg.  
Välj färg via färgdialog  
Lysfärg  
Här väljer du en lysfärg.  
Välj färg via färgdialog  
Spegelglans  
I det här området ger du objektet en spegelglans.  
Färg  
I den här listrutan väljer du spegelglansens färg.  
Välj färg via färgdialog  
Intensitet  
I detta rotationsfält kan Du definiera spegelglansens styrka i procent.  
Fördelning  
Den här funktionen används för att fördela objekt, d.v.s. för att få jämn justering.  
Du kan öppna dialogrutan om du har markerat minst tre objekt samtidigt i %PRODUCTNAME Draw eller %PRODUCTNAME Impress.  
De markerade objekten fördelas så att deras kanter eller mittpunkter ligger på samma avstånd från varandra.  
De två objekt som ligger längst från varandra, horisontellt eller vertikalt, används som fasta referenspunkter.  
De övriga objekt, som ligger mellan de yttre objekten, kan flyttas med den här funktionen.  
Horisontell  
Här definierar du avståndens horisontella fördelning.  
Ingen  
Objekten fördelas inte.  
Vänster  
Objekten placeras på jämnt avstånd från varandra räknat från objektens vänstra kant.  
Mitten  
Objekten placeras på jämnt avstånd från varandra räknat från objektens centrum.  
Avstånd  
Objekten fördelas så att alla ligger på samma avstånd från varandra.  
Höger  
Objekten placeras på jämnt avstånd från varandra räknat från objektens högra kant.  
Vertikal  
Här definierar du avståndens vertikala fördelning.  
Ingen  
Objekten fördelas inte.  
Uppe  
Objekten placeras på jämnt avstånd från varandra räknat från objektens överkant.  
Mitten  
Objekten placeras på jämnt avstånd från varandra räknat från objektens centrum.  
Avstånd  
Objekten fördelas så att alla ligger på samma avstånd från varandra.  
Nere  
Objekten placeras på jämnt avstånd från varandra räknat från objektens underkant.  
Text  
Här tilldelar du ett textritobjekt egenskaper.  
Menykommandot Text syns bara när du har skapat ett textritobjekt med hjälp av ritfunktionen.  
Rättstavning  
Med den här funktionen startar du rättstavningskontrollen. %PRODUCTNAME kan genomföra en rättstavningskontroll för ett markerat textavsnitt, aktuellt dokument, för sidhuvuden och sidfötter liksom kataloger och fotnoter.  
Rättstavningskontrollen börjar vid markörens position och fortsätter till dokumentets slut.  
En förloppsindikator visar hur kontrollen fortskrider.  
När dokumentet är slut får du en fråga om kontrollen ska fortsätta i början av dokumentet.  
Rättstavningskontrollen jämför ord för ord med posterna i ordboken.  
När skrivsättet skiljer sig åt eller om ordet inte finns i ordboken markeras ordet och dialogrutan Rättstavning visas.  
Okända men rätt stavade ord kan du lägga in i egna ordböcker.  
Original  
I dialogens huvud visas det ord som rättstavningskontrollen inte har godkänt.  
Har Du ändrat ett påträffat ord i textfältet Ord och ersatt det med ett av orden i listrutan Förslag, men vill nu ha tillbaka det "gamla" ordet?  
Då klickar Du bara på texten på raden Original så visas det "gamla" ordet där igen.  
Du kan också använda tangentkombinationen Option Alt +O.  
Ord  
Här skriver Du in den rätta stavningen av ordet som fått en anmärkning eller så väljer Du ut den rätta stavningen från listrutan Förslag.  
Som visuell hjälp visas en röd symbol med ett kryss när ordet är felaktigt i inmatningsfältet.  
Registreras ordet som riktigt visas på samma ställe en grön symbol med en bock.  
Under inmatningen visas ingen symbol.  
Kontrollera ord  
Klicka på den här kommandoknappen för att kontrollera det ändrade ordet på nytt.  
När det finns förslag för ett ändrat ord visas dessa i listrutan Förslag.  
Kontrollera ord  
Förslag  
I den här listrutan får du förslag till rätt stavning.  
Språk  
Här definierar du vilket språk som ska användas för rättstavningskontrollen av det här ordet.  
Om du ändrar språket under kontrollen så kontrolleras ordet som identifierats som felaktigt genast på det nya språket.  
Det valda språket tilldelas ordet som ett direkt teckenattribut.  
I setup-programmet kan du installera fler språkmoduler eller ta bort språkmoduler från installationen.  
Ordbok  
Här väljer du en användarordlista där du vill lägga till ordet.  
Det finns mer information om användarordlistor i dialogrutan Lingvistik.  
AutoKorrigering  
Om du klickar här läggs kombinationen av felaktigt ord och rättat ord till i AutoKorrigeringslistan.  
Mer information om AutoKorrigering.  
Synonymordlista  
Med den här kommandoknappen öppnas dialogen Synonymordlista.  
Alternativ  
Med den här kommandoknappen kommer du till dialogen Lingvistik.  
Lägg till  
Om du klickar här läggs det aktuella ordet till i den valda användarordlistan.  
Ignorera  
Genom att välja kommandoknappen Ignorera korrigeras inte det ord som stavningskontrollen har reagerat på och programmet fortsätter rättstavningskontrollen.  
Ignorera alltid  
Klicka här så korrigeras inte det ord som stavningskontrollen har reagerat på.  
Förekommer ordet på fler ställen i texten förbigås det automatiskt utan någon fråga.  
Ersätt  
Genom att välja kommandoknappen Ersätt ersätts det felaktiga ordet med det ord som Du har skrivit in direkt eller valt ut i listrutan.  
Ersätt alltid  
Klicka här när det felaktiga ordet ska ersättas med det som Du har skrivit eller valt ut.  
Förekommer ordet flera gånger i dokumentet ersätts det automatiskt utan någon fråga.  
Bakåt  
Markera kryssrutan Bakåt, när sökningen ska fortsätta från textmarkörens position i riktning mot dokumentets början.  
Statusrad  
I dialogens nedre del visas orsaken till avbrottet i den pågående rättstavningskontrollen.  
Lingvistik  
Här väljer du alternativ för rättstavningskontrollen.  
Synonymordlista  
Det är en ordlista med synonymer och du kan använda den för att söka efter ord som har samma betydelse som ett annat ord.  
Synonymordlistan stöder för tillfället inte alla språk.  
Variationer  
I detta område hittar Du urvalet med ett ord ur synonymordboken.  
Ord  
Vilket ord som visas beror på vilken position markören har när dialogrutan öppnas.  
Om synonymordlistan öppnas och markören befinner sig mitt i ett ord eller direkt framför eller bakom ett ord, så används detta ord som standard för ordsökningen.  
Betydelse  
Här får Du en lista över ett ords betydelser.  
För flertydiga ord väljer Du här den önskade betydelsen.  
Ersätt  
Här kan Du skriva in det begrepp som ska ersätta ordet, eller så kan Du överta ett ord från listrutan Synonym.  
Synonym  
Här listas de hittade liktydiga begreppen.  
Markera det önskade ersättningsbegreppet som, efter det att Du har gjort Ditt val, visas i fältet Ersätt.  
Sök  
Om de förslag som listas under Synonym inte motsvarar Dina önskemål, markerar Du den post, som bäst motsvarar det sökta begreppet, och väljer Sök.  
Det markerade begreppet används nu som utgångspunkt för sökningen efter liktydiga ord.  
Språk...  
Med den här kommandoknappen öppnar Du dialogrutan Välj språk.  
Här kan Du definiera, på vilket språk Din synonymordlista ska arbeta.  
Urval  
Här hittar Du listrutan Urval, där de tillgängliga språken listas.  
Pipett  
Med det här kommandot öppnar du fönstret Pipett med vars hjälp du kan "suga upp" färger och ersätta dem med andra färger i bitmappar och metafilsgrafikobjekt.  
När du har valt pipettverktyget kan du välja upp till fyra olika färger från ett valfritt grafikobjekt.  
De letas sedan upp i den markerade bitmappen eller metafilsgrafikobjektet och byts ut mot de färger som du har valt till höger om de sökta färgerna.  
För att du ska kunna söka och ersätta likartade färgnyanser har pipettfönstret en toleransfunktion.  
Färgtoleransen anges i procent.  
Pipett  
Växla till pipettläge genom att klicka på pipettikonen.  
När Du har klickat på ett objekt i dokumentet registreras den färg som pipettmarkören befinner sig över.  
Pipett  
Om pipettläget är aktiverat visas här den aktuella färgen som pipetten befinner sig över.  
Ersätt  
Här kan Du starta färgersättningen.  
Färgerna i en markerad bitmapp eller metafil ersätts.  
Om inga grafikobjekt av de här typerna är markerade är knappen inte tillgänglig.  
Färger  
Här kan Du definiera källfärg, tolerans och vilken färg som källfärgen ska ersättas med.  
Källfärg  
I den här kryssrutan anger Du om den visade färgen ska ersättas eller inte.  
Källfärg  
Här visas den källfärg som Du har valt.  
Tolerans  
Här kan Du ange ersättningens färgtolerans i procent.  
Ersätt med...  
Här visas en lista över alla tillgängliga färger som Du kan använda i stället för källfärgen.  
Transparens  
Om grafikobjektet redan innehåller transparenta (genomskinliga) delar kan Du välja bort transparens här.  
Transparens  
I den här listrutan väljer Du den färg som ska användas istället för transparens.  
AutoKorrigering  
I dialogrutan AutoKorrigering kan du anpassa den automatiska korrigeringsfunktionen efter dina behov.  
Du kan också låta bokstavskombinationer som Du själv anger bytas ut mot hela ord eller fraser (vilket innebär ett slags automatisk infogning av AutoText -avsnitt).  
Inställningarna av AutoKorrigeringen aktiveras när Du har skrivit färdigt teckenföljden och trycker på blankstegstangenten eller på annat sätt anger att ordet är slut.  
Varje sådan inmatning kan Du även ångra och sedan omedelbart fortsätta att skriva.  
För textdokument gäller följande: du sätter på eller stänger av den automatiska AutoKorrigeringen genom att markera respektive avmarkera menykommandot Format - AutoFormat - Under inmatningen.  
När det gäller tabelldokument hittar du motsvarande kommando under Verktyg - Cellinnehåll - AutoInmatning.  
Dessutom kan du när som helst formatera ett helt textdokument automatiskt med kommandot Format - AutoFormat - Använd.  
Info: i tabelldokument är förutom AutoKorrigeringen även AutoInmatning tillgänglig.  
Ytterligare regler för AutoKorrigering  
Någon automatisk redigering i efterhand av dokumenten är inte möjlig.  
Alternativ  
Under den här fliken definierar du de olika alternativen för AutoKorrigeringen.  
I textdokument har du tillgång till fler alternativ än i andra dokument.  
Alternativen kan användas under efterbearbetningen [E] och / eller under inmatningen [I].  
Markera motsvarande kryssrutor i kolumnerna [E] och [I].  
Om någonting t.ex. bara ska ersättas vid inmatningen, men inte vid en senare redigering av dokumentet med kommandot Format - AutoFormat - Använd, markerar du rutan i kolumnen [I] på den aktuella raden och lämnar rutan i kolumnen [E] tom.  
Markera rutorna framför samtliga rader vars alternativ programmet ska ta hänsyn till vid AutoKorrigeringen.  
Använd ersättningstabell  
Om den senast inmatade bokstavskombinationen motsvarar en förkortning i ersättningstabellen, ersätts den av motsvarande text i ersättningstabellen.  
KOrrigera två versaler i BÖrjan av ordet  
Skrivfel som "ORd" korrigeras automatiskt till "Ord ".  
Börja varje mening med stor bokstav  
Texten korrigeras på så sätt att varje ord efter slutet på en mening (representerat av t ex punkt, utropstecken, frågetecken) börjar med stor bokstav.  
Detta händer inte efter ord som består av högst två bokstäver och som följs av punkt, tankstreck, vanlig parentes eller vinkelparentes (>).  
På så sätt blir t ex a) inte oavsiktligt till A).  
Automatisk *fet* och _understruken_  
Markera den här rutan om du automatiskt vill tilldela textattributen fet och understruken.  
Skriv tecknet (_) före och efter den text som ska vara understruken.  
Tecknen själva tas bort.  
Känn igen URL  
Om detta fält är markerat försöker %PRODUCTNAME identifiera sådana teckenföljder i dokumentet som skulle kunna vara en URL.  
Varje teckenföljd som identifieras som en URL omvandlas automatiskt till en hyperlänk till denna URL.  
Mer information  
Ersätt 1 / 2... med ½...  
När Du markerar denna kryssruta byts sådana teckenkombinationer för vilka det finns en ett speciellt tecken ut mot detta tecken (exempelvis ersätts 1 / 2, 1 / 4 och 3 / 4 med ½, ¼ respektive ¾).  
Ersätt tankstreck  
Markera det här fältet om du vill göra minustecken till tankstreck.  
En teckensträng som "x[ett blanksteg][minus][ett blanksteg]xx" ersätts med "x[ett blanksteg][tankstreck][blanksteg]xx ".  
En teckensträng som "x[ett blanksteg][två minustecken]x" ersätts med "x[ett blanksteg][tankstreck]x ".  
Radera mellanslag och tabbar i början och slutet av stycke  
Om du markerar de här rutorna tas mellanslag och tabbar i början och slutet av stycken bort automatiskt.  
Radera mellanslag och tabbar mellan slutet och början på rad  
Om du markerar de här rutorna tas mellanslag och tabbar mellan början och slutet på rader bort automatiskt.  
Ersätt engelska ordningstal 1st... med 1^st...  
Om Du vill använda dig av de ordningstal som är vanliga inom engelskan, där siffrans ändelse skrivs upphöjt, markerar Du denna kryssruta.  
Övriga siffror följs av th (fourth osv).  
Ignorera dubbla blanksteg  
Om Du markerar denna kryssruta drar autokorrigeringen samman flera blanksteg till ett enda blanksteg.  
Om Du i undantagsfall i alla fall vill skriva flera blanksteg kan Du infoga ett blanksteg framför ett annat blanksteg och sedan upprepa denna procedur så ofta Du vill.  
Använd numrering  
Markera den här rutan om du vill använda en automatisk numrering eller punktuppställning vid inmatningen.  
Rader som börjar med en numrering exempelvis i form av "1 .", fortsätter i det här exemplet med "2" när Du har tryckt på returtangenten.  
Rader som börjar med ett minustecken följt av ett mellanslag eller en tabulator, blir till uppräkningar med ett bullettecken som liknar ett minustecken när Du har tryckt på returtangenten.  
Rader som börjar med ett plustecken eller en stjärna följt av ett mellanslag eller en tabulator, får ett bullettecken som Du kan välja ut när Du har klickat på kommandoknappen Redigera....  
Du korrigerar en enstaka oönskad numrering genom att trycka på Retur.  
Den automatiska numreringen aktiveras bara i stycken som formaterats med någon av styckeformatmallarna "Standard", "Brödtext" eller "Brödtext indrag ".  
Använd inramning  
Om du vill utnyttja möjligheten att skapa ett understreck automatiskt under inmatningen klickar du här.  
Understrecket skapas i form av en inramning av det föregående stycket och kan därför redigeras och raderas i det föregående styckets dialogruta Format - Stycke.  
Här följer en lista som förklarar funktionen hos de tillgängliga tecknen:  
-- -  
0,5pt Enkellinje nere  
___  
1,0pt Enkellinje nere  
===  
1,1pt Dubbellinje nere  
***  
4,5pt Dubbellinje nere  
~~~  
6,0pt Dubbellinje nere  
###  
9,0pt Dubbellinje nere  
Skriv in de tre tecknen på en tom rad och tryck sedan på returtangenten.  
Tecknen omvandlas till en inramning av det föregående stycket.  
Skapa tabell  
Med hjälp av funktionen Skapa tabell kan du infoga en tabell med några få tangenttryckningar.  
+-tecknet fungerar som kolumnavgränsare.  
Kolumnbredden definieras med minustecknet eller understrecket (_) som platshållare.  
Du kan också trycka på tabbtangenten om tabellcellen ska vara lika bred som en tabb.  
Skriv t ex följande rad i ett stycke:  
+---------------- -+-------------- -+----- - +  
Du kan direkt börja skriva text i den första cellen.  
Använd mallar  
Om autokorrigeringsfunktionen ska använda vissa styckeformatmallar automatiskt markerar du den här rutan.  
De båda tomma raderna tas bort.  
Om en sådan rad börjar med en eller flera tabulatorer får den en styckeformatmall för en underordnad rubrik motsvarande antalet tabbar.  
Ta bort tomma stycken  
Klicka här om du vill ta bort tomma stycken ur dokumentet.  
Ersätt användardefinierade formatmallar  
De användardefinierade formatmallar som används i dokumentet ersätts med fördefinierade formatmallar för textdokument.  
Den automatiska numreringen aktiveras bara i stycken som formaterats med någon av styckeformatmallarna "Standard", "Brödtext" eller "Brödtext indrag ".  
Ersätt punkttecken med  
Stycken som inleds med ett bindestreck (- minustecken), plustecken (+) eller en stjärna (*), följt av ett mellanslag eller en tabulator ersätts med bullettecknet som visas i dialogen när Du använder AutoFormat i efterhand.  
Klicka på kommandoknappen Redigera... och välj ett annat bullettecken i dialogrutan Specialtecken.  
För information om automatisk ersättning under inmatning, se Använd numrering.  
Den automatiska numreringen aktiveras bara i stycken som formaterats med någon av styckeformatmallarna "Standard", "Brödtext" eller "Brödtext indrag ".  
Ersätt raka citationstecken med typografiska  
Du kan själv ange vilka tecken som ska användas som typografiska anföringstecken genom att klicka på respektive kommandoknapp på fliken Typografiska anföringstecken.  
Kombinera enradiga stycken längre än...  
Med detta alternativ kombineras enradiga stycken som står under varandra och har formatet "Standard" till ett stycke.  
Så snart ett stycke är kortare än det inställda värdet (standardvärdet är 50% av den maximalt möjliga radlängden på sidan) kombineras det inte med det därpå följande stycket.  
Flerradiga stycken kombineras generellt sett inte ihop.  
Dialogrutan Kombinera öppnas, i vilken Du då kan ange ett större värde.  
Redigera...  
Här öppnar du en dialogruta där du kan ändra inställningarna för vald AutoKorrigering.  
Ersättning  
Här definierar du olika förkortningar för ersättning.  
Ersättningstabell  
Med posterna i ersättningstabellen definierar Du att vissa bokstavskombinationer ska ersättas med andra.  
Du kan t ex låta programmet automatiskt rätta till sådana skrivfel som Du ofta gör.  
AutoKorrigeringen kan också komma ihåg tecknens formatering.  
Om du alltid vill ha en viss text formaterad med ett visst teckensnitt formaterar du den i ett dokument med det önskade teckensnittet, markerar den sedan och öppnar dialogrutan AutoKorrigering.  
Markera inte fältet Endast text.  
I AutoKorrigering kan du ta med ramar, grafik och OLE-objekt, som är integrerade som tecken i texten.  
Välj förankringsalternativet Som tecken.  
Markera den text som står före ramen, inklusive ramen och den text som står efter ramen.  
Välj kommandot Verktyg - AutoKorrigering / AutoFormat.  
Under fliken Ersättning har den markerade texten redan infogats i fältet Ersätt.  
Skriv en förkortning och stäng dialogrutan med OK.  
Om du senare skriver förkortning i texten och trycker på mellanslagstangenten ersätter AutoKorrigering förkortningen med ersättningstexten, inklusive ram / grafik / OLE-objekt.  
För att ersättningstabellen ska kunna användas när Du skriver texten måste två villkor vara uppfyllda:  
Under Verktyg - AutoKorrigering / AutoFormat ska alternativet Använd ersättningstabell på fliken Alternativ vara markerat.  
Under Format - AutoFormat ska Under inmatningen vara markerat.  
En del ord kompletteras automatiskt även om de inte finns med i ersättningstabellen.  
Det gäller bland annat namn på veckodagar och månader.  
Om du inte vill ha den ersättningen stänger du av Komplettera ord under fliken Ordkomplettering.  
Ersätt  
Skriv här den bokstavskombination som ska ersättas automatiskt.  
med:  
Skriv här in den följd av ord, det ord eller tecken som du vill ha istället.  
Endast text  
Ersättningstexten övertar alltså den ersatta textens formatering.  
Nytt  
Med denna funktion infogas den inmatade kombinationen av ord och ersättningsord i listan.  
Knappen heter Ersätt om ordet redan finns.  
Du kan då ersätta den gamla definitionen med den nya.  
Undantag  
Här definierar du de undantag när AutoKorrigering inte ska göra några ändringar i texten.  
Definitionerna är språkberoende.  
För varje tillgängligt språk kan du definiera specifika undantag.  
Ersättning och undantag för språk:  
I listrutan väljer du det språk för vilket ersättningsreglerna / undantagen ska gälla. %PRODUCTNAME letar till att börja med efter undantag för det språk som gäller vid infogningspositionen i dokumentet.  
Därefter letar programmet igenom definitionerna för alla andra språk.  
Om du t.ex. har angett amerikansk engelska vid infogningspositionen genomförs kontrollen av ersättningsreglerna / undantagen i ordningsföljden Engelska (US) - Engelska (UK) - Alla språk.  
Förkortningar, efter vilka inga versaler följer.  
I textfältet anger Du ett ord eller en förkortning av ett ord efter vilket det kan skrivas en förkortningspunkt i texten.  
Den nästföljande bokstaven efter ett ord i en undantagslista omvandlas inte automatiskt till en stor bokstav.  
Typiska exempel i en sådan undantagslista är "etc." eller "osv. "  
Skriv också in förkortningspunkten och klicka sedan på Nytt.  
Samtliga definierade förkortningar finns med i listrutan.  
Med Radera raderar Du den aktuella förkortningen ur listan.  
Ord som börjar med två stora versaler  
Dessa ord ska alltså inte automatiskt omvandlas till ord med bara en stor bokstav av AutoKorrigeringen.  
Typiska exempel är "PC" eller "CD ".  
Alla ord som får börja med två stora bokstäver finns med i listrutan.  
Med Radera raderar du det för tillfället markerade ordet i listan.  
Nytt  
Infoga det nya undantaget i listan genom att klicka på Nytt.  
Listan sparas automatiskt och laddas automatiskt när %PRODUCTNAME startas.  
Lägg till automatiskt  
Markera den här rutan om du vill att förkortningar, som inte ska följas av stor bokstav, och ord, som börjar med två stora bokstäver, ska läggas till automatiskt i respektive lista.  
Förutsättningen för att de ska läggas till automatiskt är att alternativen KOrrigera två versaler i BÖrjan av ordet respektive Börja varje mening med en versal markerats i kolumnen [E] under Verktyg - AutoKorrigering / AutoFormat - Alternativ.  
Så snart du ändrar en korrigering som programmet gjort (t.ex. med Kommando Ctrl +Z) förs ändringen automatiskt in i respektive undantagslista. (Den här funktionen är inte tillgänglig i %PRODUCTNAME Calc.)  
Typografiska anföringstecken  
Under den här fliken definierar du utseendet för typografiska anföringstecken.  
Enkla / dubbla anföringstecken  
Här väljer Du det specialtecken på som Du vill använda för enkla och dubbla anföringstecken.  
Ersätt  
Markera den här kryssrutan om Du vill ersätta anföringstecknen.  
Datoranföringstecken ersätts med typografiska anföringstecken.  
Du kan ställa in tecknen för de typografiska anföringstecknen genom att klicka på kommandoknapparna för alternativen Vid ordets början, Vid ordets slut, Enkelt / Dubbelt anföringstecken.  
Då öppnas en dialogruta som liknar dialogrutan Specialtecken, där Du kan klicka på önskat tecken och bekräfta med OK.  
Det specialtecken som används visas bredvid kommandoknappen.  
Enkla anföringstecken används för citat inuti citat.  
Vid ordets början...  
Öppnar dialogrutan Specialtecken, i vilken Du definierar tecken vid ordets början.  
Vid ordets slut...  
Öppnar dialogrutan Specialtecken, i vilken Du definierar tecken vid ordets slut.  
Standard  
Klicka på den här kommandoknappen för att återställa tecknen vid ordets början och vid ordets slut till standardinställningen (typografiska anföringstecken).  
Snabbmenyn AutoKorrigering  
Den här snabbmenyn öppnar du genom att högerklicka på ett ord som är markerat som fel.  
<Korrigeringsförslag>  
Här visas programmets förslag till korrigering av ordet som är markerat som fel.  
Klicka på det riktiga ordet i listan.  
Rättstavning  
Med det här kommandot öppnar du dialogrutan Rättstavning.  
Lägg till  
Med det här kommandot lägger du till det markerade ordet i en av användarordlistorna.  
Ignorera alla  
Med det här kommandot raderas den röda linjen, som felmarkerar ordet, för det här ordet i hela dokumentet.  
AutoKorrigering  
Med det här kommandot visar du en undermeny med korrigeringsförslag.  
Klicka på förslaget som du vill använda så korrigeras ordet och läggs in i ersättningstabellen.  
Du kan även öppna och redigera ersättningstabellen via Verktyg - AutoKorrigering / AutoFormat - Ersättning.  
Ordet är <språkets namn>  
Det här området visas bara när flera språk är installerade och %PRODUCTNAME föreslår att ordet tillhör ett annat språk.  
Ordet kan tilldelas posten för ett annat språk.  
Stycket är <språkets namn>  
Det här kommandot visas bara när flera språk är installerade.  
Med det här kommandot kan du tilldela det andra språket ett helt stycke.  
Ordkomplettering  
Här ställer du in hur den automatiska ordkompletteringen ska fungera.  
Automatisk ordkomplettering  
Här ställer du in om du vill använda automatisk ordkomplettering och fr.o.m. vilken ordlängd den ska vara aktiv.  
Du anger ett värde vardera för minimilängd och maximalt antal ord som tas med.  
Ord som är kortare än minimal ordlängd tas aldrig med.  
Alla tillräckligt långa ord i alla dokument som du öppnat sedan du senast startade %PRODUCTNAME tas med, upp till det maximala antalet ord.  
När du börjar skriva in ett ord på nytt känner %PRODUCTNAME igen det och kompletterar det.  
Om du var på väg att skriva ett annat ord ignorerar du bara förslaget och fortsätter att skriva.  
Om du vill acceptera förslaget måste du bekräfta det med någon av tangenterna Retur, Mellanslag, Högerpil eller End.  
Sedan kan du skriva nästa ord. (I fältet Acceptera med väljer du med vilken tangent du vill bekräfta).  
Eftersom ordkomplettering sker fr.o.m. den tredje bokstaven som du skriver visas inte alltid det önskade ordet med en gång.  
Om det finns flera ord i AutoKorrigeringens minne som börjar med samma bokstäver kan du titta på alternativen och välja ett av dem.  
När ordkompletteringen visas, trycker du på Kommando Ctrl +Tabb.  
Ett nytt förslag visas direkt.  
Detta sker tills det inte finns några fler förslag.  
Med Kommando Ctrl +Skift+Tabb bläddrar du genom förslagen åt andra hållet.  
Därför kan det ta en stund innan %PRODUCTNAME hinner sammanställa en aktuell lista i bakgrunden om texterna är långa.  
Listan raderas när du avslutar %PRODUCTNAME.  
Visa förslag  
Om den här rutan är markerad visas förslagen från den automatiska ordkompletteringen antingen som markerad text eller som tipshjälp när du skriver in text.  
Samla förslag  
När det här alternativet är markerat samlas förslagen i en redigerbar lista som visas i listrutan på den här fliken.  
Oändliga förslag  
Efter det sista förslaget visas det första igen osv.  
Om alternativet inte är markerat kan Du inte bläddra kontinuerligt utan bara till första och sista förslaget.  
Tillfoga mellanslag  
När det här alternativet är markerat infogas ett blanksteg efter en automatisk ordkomplettering.  
Visa som tipshjälp  
Om det här alternativet är markerat visas förslagen från den automatiska ordkompletteringen endast som tipshjälp.  
Min. ordlängd  
I det här rotationsfältet anger du värdet för minsta ordlängd för de ord som ska sparas.  
Max poster  
I det här rotationsfältet kan du definiera hur många ord som maximalt ska sparas.  
Acceptera med  
Här kan Du välja vilken tangent Du ska acceptera det aktuella förslaget från den automatiska ordkompletteringen med  
Ordlista  
Listan bibehålls tills %PRODUCTNAME stängs.  
Du kan markera ord i listan genom att klicka på dem eller avmarkera enskilda ord.  
Om Du klickar på ett ord och samtidigt trycker ned skifttangenten markeras alla ord mellan det senast markerade ordet och det ord som Du klickar på.  
Du kan kopiera alla markerade ord i listan till urklippet med Kommandot Ctrl +C.  
Från urklippet kan du sedan klistra in orden i t.ex. ett textdokument och spara det som en referensordlista.  
Textdokumentet kan du vid behov utöka eller redigera manuellt.  
Om Du vid ett senare tillfälle ska skriva en text i %PRODUCTNAME och behöver de sammanställda orden igen, kan Du markera alternativet Samla förslag på fliken Ordkomplettering och sedan öppna referensordlistan.  
Dina ord kommer då med i listan.  
Avmarkera sedan alternativet Samla förslag igen och växla till det nya textdokumentet som Du ska skriva.  
När Du skriver har Du tillgång till förslag från referensordlistan.  
Om den automatiska rättstavningskontrollen är aktiverad samlas bara ord som rättstavningskontrollen känner igen.  
Radera post  
Om du klickar på den här kommandoknappen tas alla ord som är markerade i ordlistan bort.  
Numrering / punktuppställning  
Med den här funktionen kan du infoga numreringar eller punktuppställningar i ett dokument.  
I %PRODUCTNAME Impress kan du använda automatisk numrering för en - eller flerradiga stycken.  
För dispositionsobjekt (Stylist) kan upp till nio numreringsnivåer användas, för textobjekt upp till tio.  
Den tilldelade numreringen uppdateras automatiskt efter ändringar i de numrerade styckena.  
I %PRODUCTNAME Draw kan du använda automatisk numrering för en - eller flerradiga stycken.  
För dispositionsobjekt (Stylist) kan upp till nio numreringsnivåer användas, för textobjekt upp till tio.  
Den tilldelade numreringen uppdateras automatiskt vid ändringar i de numrerade styckena.  
I %PRODUCTNAME Writer kan du använda automatisk numrering för en - eller flerradiga stycken.  
Numreringen kan göras i efterhand eller medan texten skrivs. %PRODUCTNAME Writer stöder upp till tio numreringsnivåer.  
Den tilldelade numreringen uppdateras automatiskt efter ändringar i de numrerade styckena.  
Det går även att infoga stycken utan numrering och att via tangentbordsinmatningar undanta enstaka stycken från löpande numrering, så att en nivå kan bestå av flera stycken.  
Markera de stycken som numreringen eller punktuppställningen ska gälla för.  
Om inga särskilda stycken markerats gäller ändringen för aktuellt stycke.  
Öppna dialogrutan och välj en punkt, en numreringstyp, en disposition eller ett grafikobjekt för visningstypen uppställning eller numrering.  
Om du inte anger något val utan avslutar dialogrutan med OK numreras det aktuella stycket med dialogrutans förinställningar.  
Då stängs även dialogrutan.  
Du kan lägga till fler dispositionsnivåer genom att ställa markören på en nivå direkt efter punktuppställningstecknet och trycka på tabbtangenten.  
Om markören står i en dispositionsnivå utan att något tecken eller ord är markerat, gäller ändringarna som du gör i dialogrutan Numrering / punktuppställning för en hel nivå.  
Om däremot minst ett tecken är markerat, gäller en ändring bara för det aktuella stycket.  
Ändringar som du gör i dialogrutan Numrering / punktuppställning gäller, oavsett dispositionsnivå, bara för det aktuella stycket.  
När markören står i en numrering eller punktuppställning visas ikonerna för redigering av numreringen eller punktuppställningen på numreringsobjektlisten objektlisten objektlisten.  
Med ikonen Redigera numrering Punktuppställningstecken öppnar du dialogrutan Numrering / punktuppställning, där du kan definiera eller ändra egenskaperna för en numrering eller punktuppställning.  
I dialogrutan Numrering / punktuppställning finns följande flikar.  
Radera  
Med det här alternativet tar du bort automatisk numrering / punktuppställning i det aktuella stycket eller i de markerade styckena.  
Den här funktionen är även tillgänglig via ikonen på objektlisten.  
Punkter  
Här kan du välja en speciell punkt.  
Du kan göra fler inställningar under flikarna Position (respektive Indrag och avstånd för presentationsobjektmallar) och Alternativ.  
Punkterna är identiska med de grafikobjekt som finns i temat Punkter i Gallery.  
Om du lägger till fler grafikobjekt i temat Punkter i Gallery visas även dessa i den här dialogrutan.  
Urval  
Här väljer du önskad punkt.  
Numreringstyp  
Här kan du välja önskad numreringstyp.  
Du kan göra fler inställningar under flikarna Position (respektive Indrag och avstånd för presentationsobjektmallar) och Alternativ.  
Urval  
Välj önskad numreringstyp här.  
Disposition  
Här kan du bestämma dispositionstyp för en numrering / punktuppställning med flera nivåer.  
Urval  
Välj önskad disposition här.  
Grafik  
Här kan du välja grafik som tecken för en punktuppställning..  
Du kan göra fler inställningar under flikarna Position (resp. Indrag och avstånd för presentationsobjektmallar)  
Urval  
Välj ett grafikobjekt här.  
Länka grafik  
Markera den här rutan om du vill länka ett grafikobjekt till dokumentet.  
Om rutan inte är markerad, integreras grafikobjektet i dokumentet.  
Det är bättre än att länka om dokumentet öppnas på en dator där Gallery inte är tillgängligt.  
Alternativ  
Här definierar du visningstyp för numreringar och punktuppställningar.  
Du kan definiera formateringar för varje dispositionsnivå för sig eller för alla nivåer samtidigt.  
Nivå  
Denna listruta används för att välja en dispositionsnivå, för vilken Du sedan kan ställa in alternativ i området Format.  
Aktuell formatering visas i förhandsvisningsfältet.  
Om Du väljer alternativ "1 -10" kan Du ange inställningar för alla nivåer samtidigt.  
Format  
I detta område definierar Du början för och typen av numrering för den eller de valda nivåerna.  
Numrering  
I detta kombinationsfält väljer Du numreringstyp för den eller de aktuella nivåerna.  
Urval  
Funktion  
1, 2, 3,...  
Arabiska siffror  
A, B, C,...  
Versaler  
a, b, c,...  
Gemener  
I, II, III,...  
Versala romerska siffror  
i, ii, iii,...  
Gemena romerska siffror  
A,...  
AA,...  
AAA,...  
Antalet bokstäver anger dispositionsnivån.  
Andra numreringen på tredje nivån blir alltså "BBB".  
a,... aa,... aaa,...  
Antalet bokstäver anger dispositionsnivån.  
Tredje numreringen på andra nivån blir alltså "cc".  
Punkt  
Ett specialtecken (punkt) placeras före första raden i stycket.  
Om du väljer den här typen kan du öppna dialogrutan Specialtecken via kommandoknappen... och välja en punkt.  
Punkternas storlek anpassas till radhöjden om du inte själv har definierat en teckenformatmall med egen teckenstorlek för punkter.  
Grafik  
Grafiken kan definieras via kommandoknappen Urval....  
Grafik länkad  
Om du vill infoga ett grafikobjekt, som du använder för en punktuppställning / numrering, som en länk i dokumentet markerar du det här alternativet.  
Något länkat grafikobjekt är då inte tillgängligt.  
Ingen  
Inga numreringstecken.  
Bara tecken som definierats som avgränsare visas vid radens början.  
Formateringsmöjligheterna för en numrering eller punktuppställning varierar beroende på om du valt en siffra, en punkt eller ett grafikobjekt som tecken.  
Följande fält visas därför bara när motsvarande alternativ valts under Numrering.  
Framför  
Om vissa tecken ska placeras framför numreringen anger du dem här.  
Med "Till" erhålls numreringen "Till 1 ".  
Bakom  
Om vissa tecken ska placeras före numreringen ska dessa anges här.  
För vissa numreringstyper placeras som standard en punkt mellan numreringstecknet och radens början.  
Denna standard kan Du skriva över eller utöka.  
Med ".)" erhålls numreringen "1.) ".  
Teckenformatmall  
I det här kombinationsfältet kan du välja en teckenformatmall för numreringen om du vill.  
Du kan t.ex. även välja mer ovanliga teckenuppsättningar.  
Fullständig  
I detta rotationsfält kan Du ange hur många överordnade nivåer som ska visas för den eller de aktuella numreringsnivåerna.  
Om Du t ex ställer in värdet 2 för den tredje nivån erhålls en numrering typ "1.1." för denna nivå.  
Det värde som kan ställas in via detta rotationsfält begränsas av aktuell numreringsnivå.  
Börja med  
Här definierar du vilket nummer som numreringen ska börja med.  
Färg Färg  
Om du har valt alternativet punkt under Numrering kan du välja färg till punkten här.  
Om du har valt alternativet punkt under Numrering kan du välja punktens färg här.  
Relativ storlek Relativ storlek  
Om du har valt alternativet punkt under Numrering kan du ställa in punktens storlek här.  
Storleken anges i förhållande till aktuell teckenhöjd i stycket.  
Om du valt alternativet punkt under Numrering kan du ställa in punktens storlek här.  
Storleken anges i förhållande till aktuell teckenhöjd i stycket.  
Tecken  
Genom att klicka på kommandoknappen... öppnar du dialogrutan Specialtecken där du kan leta fram ett punkttecken.  
Den här funktionen är bara tillgänglig om du har valt alternativet punkt under Numrering.  
Om Du har valt alternativet Grafik under Numrering:  
Urval...  
När Du klickar på denna kommandoknapp kan Du välja grafik från Gallery.  
Då öppnas en undermeny där Du kan välja bland alternativen Från fil... och Gallery.  
Via posten Från fil... öppnas dialogrutan Länka där Du kan välja ett grafikobjekt.  
Denna dialogruta är upplagd på samma sätt som Infoga grafik.  
Via posten Gallery öppnas en popup-meny, där Du kan välja ett grafikobjekt direkt från Gallery.  
Bredd  
Här definierar Du grafikobjektets bredd.  
Höjd  
Här definierar Du grafikobjektets höjd.  
Synkronisering  
Om Du markerar denna kryssruta bibehålls grafikobjektets höjd - / breddförhållande vid storleksförändring.  
Justering  
Här bestämmer Du hur grafikobjektet ska justeras.  
Alla nivåer  
Här kan Du ange en fortlöpande numrering för alla nivåer.  
Fortlöpande numrering  
När Du har markerat denna kryssruta numreras alla nivåer fortlöpande.  
Position  
Här formaterar du styckena i dispositionen.  
Den här funktionen är tillgänglig för både kapitelnumreringar (Verktyg - Kapitelnumrering) och stycken som ska förses med en numrering eller punktuppställning (Format - Numrering / punktuppställning).  
Om du redigerar en kapitelnumreringar är de formateringar som du har valt under fliken Position indirekta formateringar med mallar eftersom formateringarna påverkar de styckeformatmallar som har tilldelats under fliken Numrering.  
Om du redigerar en numrering eller punktuppställning är de formateringar som du valt under fliken Position direkta formateringar som inte är bundna till en viss mall.  
Nivå  
Därefter kan Du göra inställningar på denna flik.  
Aktuell formatering visas i förhandsvisningsfältet.  
Välj alternativet "1 -10" om Du vill ange inställningar för alla nivåer samtidigt.  
Position och avstånd  
I detta område ställer Du in den exakta placeringen av dispositionsnivåtecknen och de nivåindelade styckena för varje dispositionsnivå.  
Tänk på att inställningarna som du gör här påverkar det aktuella styckets formatering, som definieras under Format - Stycke... - Indrag och avstånd för en punktuppställning / numrering.  
De inställningar som du gör här påverkar det aktuella styckets formatering, som definieras under Format - Stycke - Indrag och avstånd för en punktuppställning / numrering.  
Vid en kapitelnumrering ställer du in formateringen under motsvarande flik för styckeformatmallen.  
När du definierar värden för avståndet mellan text och textram under fliken Position kommer värdena för indrag av stycket som finns i området Indrag under fliken Indrag och avstånd att anpassas på motsvarande sätt.  
Om du sedan anger andra värden där, kommer inte längre någon hänsyn att tas till de inställningar som du har gjort här för numrering / punktuppställning.  
När Du definierar värden för avståndet mellan numreringstecknen och sidmarginalen med hjälp av Indrag på fliken Position kommer värdena för indrag av stycket som finns i området Indrag på fliken Indrag och avstånd att läggas till.  
Tidigare styrdes radindragen för stycken med hjälp av en numrering.  
I %PRODUCTNAME anpassas inställningarna i styckedialogrutan under Indrag och avstånd och i numreringsdialogrutan under Position automatiskt till respektive programversion.  
Indrag  
I detta rotationsfält definierar Du avståndet mellan det vänstra styckeindraget och vänstermarginalen för numreringstecknet.  
Om Du inte har ställt in något styckeindrag på fliken Indrag och avstånd (Från vänster = 0 cm) motsvarar indraget avståndet mellan sidans vänstermarginal och numreringstecknet.  
I det här rotationsfältet definierar du avståndet mellan den vänstra textramen och vänster styckemarginal respektive numreringstecken.  
Det här värdet fylls i som vänster styckeindrag under fliken Indrag och avstånd.  
Relativ  
Om Du har markerat detta alternativ tolkas det värde som Du har angett under Indrag relativt till den överordnade dispositionsnivån.  
För den första dispositionsnivån har detta fält ingen effekt.  
Avstånd till text  
Här ställer Du in avståndet mellan numreringstecknet och texten.  
Minimum avstånd numrering <-> text  
Här kan Du definiera ett minimiavstånd mellan numreringstecknet och texten efter detta tecken.  
Detta miniminavstånd kan t ex se till att det blir ett tillräckligt avstånd mellan numreringstecknet och texten när numreringstecknet är högerjusterat.  
Placering av numrering  
Här definierar Du dispositionsnivåtecknenas placering.  
Du väljer mellan vänsterjusterad, högerjusterad eller centrerad placering.  
Vid placeringen tas alltid hänsyn till det minimiavstånd mellan text och numrering som Du angett under Minimum avstånd numrering <-> text.  
Detta innebär att en centrerad eller högerjusterad placering bara är möjlig i den mån som detta minimiavstånd tillåter det.  
Detta placeringsalternativ hänför sig endast till numreringstecknen och inte till alla kapitelrubrikerna eller det numrerade stycket.  
Du definierar styckets placering på fliken Placering.  
Standard  
Med denna knapp återställer Du värdena för avstånd och indrag till de fördefinierade standardvärdena som finns i programmet.  
Makro  
Här administrerar och redigerar du makron.  
Makronamn  
Du kan också ange ett namn för ett nytt makro.  
I den här listrutan visas de makron som finns i den modul som du har markerat i listrutan Makro från.  
Markera ett makro om du vill redigera eller visa det.  
Makro från  
I denna listruta väljer Du ut den modul som innehåller ett makro som Du vill redigera eller som Du vill skapa ett nytt makro för.  
Om Du vill föra in ett makro i en bestämd fil måste Du först öppna filen.  
Beskrivning  
Här ser du beskrivningen av det markerade makrot, om det finns någon.  
Kör  
Genom att trycka på knappen kör Du det befintliga makrot som Du har markerat i området Makronamn.  
Tilldela  
Med den här kommandoknappen öppnar du dialogrutan Anpassa.  
Där kan du tilldela en meny, ett tangentkommando eller en händelse det nya makrot.  
Redigera  
Startar Basic-IDE och öppnar den markerade makromodulen.  
Nytt / Radera  
Raderar den för tillfället markerade posten eller används för att skapa en ny post när du skrivit in ett nytt namn.  
Den här kommandoknappen heter Nytt när du har angett ett nytt namn i textfältet Makronamn.  
Klicka på knappen om du vill ange ett nytt makro.  
Detta är förberett för dina inmatningar genom att textmarkören redan befinner sig i en subrutin (Sub / End Sub).  
Om du har markerat ett befintligt makro i listrutan Makronamn så heter den här kommandoknappen Radera.  
Makrot tas bort från källtexten.  
Administrera  
Med hjälp av dialogrutan Administrera administrerar du modulerna, dialogrutorna och biblioteken.  
Du kan aktivera och inaktivera enstaka bibliotek, lägga till eller radera befintliga bibliotek och definiera nya.  
Du kan också definiera, redigera och radera moduler och dialogrutor.  
Fliken Modul  
Här organiserar Du moduler och dialogrutor.  
Modul / Dialog  
Klicka på Ny dialog eller Ny modul.  
Därefter måste du ange ett namn för den nya modulen eller den nya dialogen.  
Modul / Dialog  
Här visas de befintliga modulerna och dialogerna i programmet och i öppnade dokument.  
Om du vill lägga till ett nytt element markerar du ett bibliotek.  
I denna listruta flyttar och kopierar Du element genom att dra och släppa dem mellan programmet och det öppnade dokumentet.  
Dra ett element till det ställe i listrutan som Du vill flytta det till.  
En linje under markören visar exakt var elementet kommer att infogas när Du släpper musknappen.  
Om Du vill kopiera håller Du ned tangenten Alternativ Alt samtidigt som Du drar.  
Redigera  
Klicka på den här kommandoknappen om du vill redigera den markerade modulen eller dialogen.  
Då visas %PRODUCTNAME Basic-gränssnittet.  
Ny modul  
Klicka här om du vill skapa en ny modul.  
Modulen fogas in i det bibliotek som markerats i listrutan.  
Du kan ange ett namn i en dialogruta.  
Du ser därefter %PRODUCTNAME Basic-gränssnittet.  
Ny dialog  
Klicka här om du vill skapa en ny dialogruta.  
Dialogrutan infogas i det bibliotek som markerats i listrutan och ges det namn som skrivits in i textfältet.  
Därefter visas %PRODUCTNAME Basic-gränssnittet.  
Fliken Bibliotek  
Här förvaltas de bibliotek i vilka moduler och dialogrutor är sammanfattade.  
Enskilda bibliotek kan aktiveras och inaktiveras, nya kan infogas och olika bibliotek kan redigeras och raderas.  
Bibliotek  
Det kan röra sig om ett program eller ett av de öppna dokumenten.  
Bibliotek  
I den stora listrutan nedanför visas namnen på biblioteken.  
Inaktivera varje enskilt bibliotek genom att avmarkera det.  
Redigera  
Klicka på den här kommandoknappen om du vill redigera det markerade biblioteket.  
Du ser därefter %PRODUCTNAME Basic-gränssnittet.  
Lösenord  
När du klickar på den här kommandoknappen kommer du till dialogrutan Ändra lösenord.  
Nytt  
Klicka här om Du vill skapa ett nytt bibliotek.  
I dialogrutan Nytt bibliotek anger Du namnet på det nya biblioteket.  
Namn  
Ange det nya bibliotekets namn.  
Skapa separata filer  
Markera detta fält om det nya biblioteket ska sparas som en fristående fil (i {installpath} / user / basic).  
Makron som sparats som separata filer laddas inte automatiskt när %PRODUCTNAME startas, utan måste aktiveras med anrop från andra makron eller "för hand".  
Lägg till  
Här väljer Du ett befintligt bibliotek som ska läggas till i listen.  
Denna dialogruta är i allt väsentligt densamma som dialogrutan Öppna.  
Välj önskat bibliotek och klicka på Öppna.  
Här kan Du ange olika alternativ.  
Ändra lösenord  
I den här dialogrutan kan du skydda ett makro med hjälp av ett lösenord.  
Du kan ange ett nytt lösenord eller ändra ett befintligt.  
Gammalt lösenord  
Här finns textfältet där det gamla lösenordet ska skrivas.  
Lösenord  
Ange det gamla lösenordet här (om du har något).  
Nytt lösenord  
I det här området definierar du det nya lösenordet.  
Lösenord  
I det här textfältet anger du det nya lösenordet.  
Bekräfta  
I det här textfältet upprepar du det nya lösenordet.  
Lägg till bibliotek  
I den här dialogrutan kan Du lägga till %PRODUCTNAME Basic-bibliotek från en i förhand vald fil till de befintliga biblioteken.  
Filnamn:  
I listrutan ser du de bibliotek som filen innehåller.  
Markera de bibliotek som du vill lägga till genom att markera rutan framför namnet.  
Alternativ  
I det här området gör Du ytterligare preciseringar.  
Infoga som referens (endast läsning)  
Markera den här rutan om de markerade biblioteken bara ska integreras för läsning.  
På det här sättet kan flera användare ha åtkomst till samma bibliotek som är placerade centralt på en företagsserver.  
Första gången ett makro körs när du har startat om %PRODUCTNAME, läses de aktuella biblioteken in av servern.  
Spara som separat fil  
Markera den här kryssrutan om en kopia av biblioteket ska sparas som separat fil på hårddisken.  
Ersätt existerande bibliotek  
Om Du markerar den här kryssrutan, ersätts befintliga bibliotek av nyinlästa som har samma namn.  
Anpassa  
Den här funktionen ger möjlighet till individuell programanpassning.  
Gränssnitten i %PRODUCTNAME är i stor utsträckning möjliga att konfigurera för olika aktiverade dokumenttyper.  
Vidare kan Du ändra tangentkombinationerna för kortkommandon och skapa nya symbollister.  
Du kan anpassa %PRODUCTNAME globalt för alla dokument av en viss dokumenttyp, men Du kan också koppla en viss konfiguration till ett valfritt %PRODUCTNAME -dokument.  
Globala anpassningar gäller för alla dokument av en och samma typ.  
Om du gör en anpassning av t.ex. symbollisterna, och det aktiva dokumentet är ett textdokument, gäller den här anpassningen fortsättningsvis när det aktiva dokumentet är ett textdokument.  
Om Du vill att en anpassning ska gälla bara för ett enskilt, speciellt dokument, kan Du lägga till konfigurationen som fil till dokumentfilen (se nedan).  
Alternativt kan du öppna dialogrutan Anpassa genom att klicka på en symbollist med höger musknapp.  
När Du laddar egendefinierade menyer, ikonlister och tangentkonfigurationer från filer, tänk då på att Du först måste byta till motsvarande flik innan Du klickar på laddningsikonen.  
Om Du t ex vill ladda en egen tangentkombination från en fil, måste Du byta till fliken Tangentbord.  
Om Du t ex vill ändra innehållet på den objektlist eller menylist som Du ser när Du har ett dokument öppet, måste Du först ladda ett textdokument innan Du redigerar listen i fråga.  
Om Du t ex har ändrat tangentkombinationerna för kortkommandon, kan Du spara denna nya tangentanvändning som en fil.  
Klicka i så fall på kommandoknappen Spara på fliken Tangentbord.  
Ange t ex Tangenter.cfg som namn.  
Senare, när Du t ex har gjort en komplett nyinstallation av %PRODUCTNAME på en ny dator, kan du åter ladda tangentkonfigurationen (kommandoknappen Ladda på fliken Tangentbord).  
I Anpassa-dialogrutan redigerar du alltid konfigurationen av den aktuella modulen (%PRODUCTNAME Writer, %PRODUCTNAME Calc och så vidare).  
Följande steg-för-steg-anvisningar hittar du i %PRODUCTNAME -hjälpen:  
Ändra en symbollist  
Ändra tilldelning av tangentkombinationer  
Ändra en meny.  
Meny  
Under den här fliken kan du anpassa menyerna efter dina personliga behov.  
Spara den nya menyindelningen med ett beskrivande namn, så att du ladda menyerna senare igen.  
Snabbmenyerna går inte att ändra.  
Menyposter  
Här visas menyposternas struktur och bredvid den de tilldelade funktionerna.  
Tilde-tecknet står framför respektive tecken som visas med en understrykning i den färdiga menyn.  
I de andra indragna nivåerna visas menyernas innehåll.  
Här redigerar Du menylisten i det aktuella sammanhanget.  
Det betyder att Du för att kunna bearbeta den menylist som är aktiv när Du arbetar med ett textdokument först måste göra ett textdokument till aktuellt dokument.  
Motsvarande gäller också när Du ska bearbeta symbollister och snabbtangenter.  
Genom att dra och släppa kan du ändra placeringen av de enskilda menyalternativen.  
Markera ett menyalternativ, håll ner musknappen och dra det till önskat ställe.  
Medan du drar med musen visar en hjälplinje var menyalternativet kommer att infogas när du släpper musknappen.  
Skapa ett nytt menykommando genom att klicka på knappen Nytt.  
En ny undermeny skapas med knappen Ny meny.  
Om du vill skapa ett menyalternativ på den översta hierarkinivån, t.ex. bredvid menyn Hjälp, måste du stänga den tidigare menyn (menyn omedelbart till vänster), markera den och sedan klicka på knappen Ny meny.  
Du öppnar och stänger menyn genom att dubbelklicka på namnet.  
Du kan ändra namnet på ett markerat menyalternativ genom att klicka på det och sedan vänta ett ögonblick.  
Nu är inte längre hela raden markerad, utan bara namnet.  
Redigera namnet på samma sätt som vid textfält.  
Om du vill tilldela ett menyalternativ en ny funktion markerar du posten i listrutan med musen och väljer sedan önskad funktion i området Funktioner.  
När du klickar på kommandoknappen Ändra övertas ändringen av menyalternativet.  
Funktioner  
Kategori  
Här kan Du välja den kategori ur vilken Du vill tilldela ett menyalternativ en funktion.  
Funktion  
Välj den funktion som Du vill tilldela ett menyalternativ.  
Den streckade linje som står som det översta alternativet i fältet Funktion, används för att foga in en underindelning i en meny.  
Nytt  
Här kan du skapa ett nytt menyalternativ.  
Klicka i listrutan Meny på det ställe där det nya kommandot ska infogas och bekräfta med Nytt.  
Ny meny  
Här kan Du skapa ett nytt menyalternativ för en undermeny.  
Istället för att bekräfta med kommandoknappen Ny väljer Du istället Ny meny.  
Ändra  
Här kan du ändra ett befintligt menyalternativ.  
Markera det menyalternativ som ska ändras, välj önskad kategori och funktion och bekräfta med Ändra.  
Uppåtpil  
Med denna knapp flyttar Du menyalternativen uppåt.  
Menyalternativen flyttas stegvis, dvs menyalternativ för menyalternativ.  
Med kommandoknappen kan Du ändra strukturen i Din menylist, genom att t ex flytta menyalternativet Rättstavning från Verktyg-menyn till Arkiv-menyn.  
Uppåtpil  
Nedåtpil  
Med den här knappen flyttar du menyalternativ nedåt.  
De flyttas stegvis.  
Varje gång du klickar på kommandoknappen flyttas det markerade menyalternativet ett steg nedåt.  
På detta sätt kan du t.ex. flytta ett menyalternativ från menyn Redigera till menyn Infoga.  
Nedåtpil  
Du kan även flytta menyalternativ till andra ställen i menystrukturen genom att dra och släppa dem.  
Ladda...  
Med denna symbol kommer Du till dialogrutan Ladda menykonfiguration.  
Denna dialogruta har en uppbyggnad som liknar dialogrutan Öppna.  
Du kan ladda en tidigare sparad menykonfiguration för fortsatt användning.  
En konfiguration gäller tills den ersätts av en ny konfiguration.  
Spara...  
Där kan du spara din personliga konfiguration.  
Tangentbord  
Under den här fliken kan du anpassa tangentbordet efter dina behov.  
Tangentkombinationer  
I den här listrutan ser Du till vänster de tangenter eller tangentkombinationer som Du kan använda till att konfigurera tangentbordet.  
Till höger om dem hittar Du inom hakparenteser tillhörande funktioner.  
Du redigerar här kortkommandona i det aktuella sammanhanget.  
Det betyder att Du för att kunna redigera de kortkommandon som Du vill använda på ett textdokument först måste göra ett textdokument till aktuellt dokument.  
Först därefter kan Du öppna dialogrutan Anpassa.  
Detsamma gäller även för redigering av symbollisterna och menyerna.  
En steg-för-steg-handledning i hur Du anpassar kortkommandon finns i beskrivningen av hur Du gör en Tilläggsfunktion till stavningskontrollen med hjälp av en tangenttryckning.  
Funktioner  
Med hjälp av listrutorna Kategori och Funktion väljer Du här en funktion som du vill tilldela en viss tangent eller tangentkombination.  
Kategori  
Den här listrutan visar vilka funktionsområden Du kan välja bland, inklusive egenprogrammerade Basic-bibliotek.  
Funktion  
I den här listrutan visas de funktioner som hör till det markerade funktionsområdet.  
Tangenter  
Om en tangentkombination redan har tilldelats den valda funktionen så visas den i det här fältet.  
Ändra  
Med den här kommandoknappen tilldelar Du den valda funktionen den tangent eller tangentkombination som Du har angett i listrutan Tangentbord.  
Om tangenten eller tangentkombinationen redan används för en annan funktion, kommer den gamla användningen automatiskt att skrivas över av den nya utan att Du behöver bekräfta detta.  
Ändringarna verkställs dock inte förrän Du stänger dialogrutan genom att klicka på OK.  
Ladda...  
Med den här kommandoknappen öppnar Du dialogrutan Ladda tangentbordskonfiguration, i vilken Du kan öppna en tidigare sparad tangentbordskonfiguration.  
Den här dialogrutan motsvarar dialogrutan Öppna.  
Spara...  
Med den här kommandoknappen öppnar du dialogrutan Spara tangentbordskonfiguration där du kan spara din personliga konfiguration.  
Statuslist  
Under den här fliken anger du vilka data som ska visas på statuslisten.  
Statuslist  
Genom att markera motsvarande kryssruta i denna stora listruta definierar Du vilken information som ska visas på statuslisten.  
Ladda...  
Den är uppbyggd på samma sätt som dialogrutan Öppna.  
Spara...  
Med den här kommandoknappen kommer du till en dialogruta där du kan spara din statuslistkonfiguration.  
Symbollister  
Här kan du konfigurera symbollisterna.  
Om Du inte ser den symbollist som ska redigeras stänger Du först dialogrutan Anpassa, laddar sedan ett lämpligt dokument eller öppnar ett nytt tomt dokument av rätt typ där Du kan se symbollisten och öppna därefter dialogrutan Anpassa på nytt.  
Synliga symbollister  
Här ser du namnen på alla huvudsymbollisterna.  
Genom att markera kryssrutorna definierar du vilka lister som ska visas.  
Om du avmarkerar en kryssruta framför en post visas inte motsvarande list mer.  
Alla symbollister som visas under fliken Symbollister har en särskilt lättanvänd snabbmeny.  
Via undermenyn Anpassa kommer du till fliken Symbollister.  
Med menypunkten Redigera öppnar du dialogrutan Redigera symbollister.  
Du kan också öppna den via Visa - Symbollister - Redigera.  
Under Synliga kommandoknappar finns en lista över alla ikoner som listen innehåller, indelad i visade och dolda ikoner.  
Synliga ikoner är markerade med en bock.  
Genom att klicka enkelt med musen på en av ikonerna i listan visas eller döljs ikonen.  
Alternativ  
Innehåll  
Här kan Du välja mellan visningssätten Ikon, Text eller Ikon+Text för symbollisterna.  
Du kan definiera en individuell inställning för varje list.  
Markera önskad list i listrutan Symbollister och välj önskat visningssätt i listrutan Innehåll.  
Ny  
Här kan du skapa nya egna symbollister.  
Redigera...  
Med kommandoknappen Redigera... öppnar du dialogrutan Redigera symbollister.  
Du drar ikoner från symbolfönstret och släpper dem på symbollisterna och kan flytta eller ta bort ikoner som redan är placerade där.  
En del av ikonerna saknar grafisk utformning.  
Där kan du välja ut ett grafikobjekt som du kan tilldela ikonen.  
Förinställning  
Genom att klicka på denna kommandoknapp återtar Du ändringarna i den list som markerats under Symbollister.  
Ladda...  
Om du klickar på den här kommandoknappen öppnas dialogrutan Ladda symbollistkonfiguration, som är uppbyggd på samma sätt som dialogrutan Öppna.  
Spara...  
Med den här kommandoknappen kommer du till en dialogruta där du kan spara din symbollistkonfiguration.  
Om Du har redigerat några symbollister och sedan klickar på Återställ, återställs omedelbart och oåterkalleligt de ändringar som Du har gjort i samtliga symbollister.  
Redigera symbollister  
Här redigerar du symbollisterna.  
Välj först ett område och en funktion i den nedre delen av dialogrutan.  
I den övre delen av dialogrutan visas då automatiskt den tillhörande kommandoknappen intryckt.  
Du måste eventuellt rulla för att se den.  
Dra den intrycka kommandoknappen från dialogrutan och släpp den på symbollisten.  
Lägg också märke till snabbmenyn på symbollisten.  
De är uppdelade efter de som för tillfället är synliga och de som inte är synliga.  
De synliga ikonerna är markerade med en bock.  
Genom att klicka med musen på en ikon utan bock blir ikonen synlig på listen.  
Ikoner  
Här finns kommandoknapparna som hör till kategorin som är markerad i listrutan Kategori.  
Varje funktion som finns i listrutan Funktion motsvarar en kommandoknapp.  
Funktioner  
Kategori  
Här markerar du den kategori som ikonen eller motsvarande funktion tillhör.  
Funktion  
Här markerar du den funktion som är definierad i kategorin som du valde innan.  
Ikoner...  
I dialogrutan kan du redigera den markerade funktionsknappen.  
Dialogrutan går bara att öppna när du har markerat en ikon eller en kommandoknapp.  
Redigera kommandoknapp  
I den här dialogrutan tilldelar du den funktionsknapp som du har markerat tidigare en valfri ikon.  
Det finns olika ikoner att välja mellan.  
Välj den ikon som du vill använda för att visa funktionsknappen och bekräfta genom att klicka på OK.  
Du måste dock kopiera dem i BMP-format till mappen "{installpath} / share / config / symbol".  
Varje gång Du startar dialogrutan Redigera kommandoknappar söks mappen automatiskt igenom efter nya ikoner med hjälp av %PRODUCTNAME.  
Storleken på ikonerna får inte överstiga 30x30 pixlar och 256 färger.  
Funktion:  
Här ser Du beskrivningen av funktionsknappen.  
Du ändrar beskrivningen genom att ange ett nytt namn.  
Standard  
När Du klickar på denna knapp kan Du ångra de ändringar som Du har gjort för de funktionsknappar som markerats under Ikoner.  
Händelser  
Makrona utförs då den valda händelsen inträffar.  
Händelse  
I listrutan Händelse väljer du ut den programhändelse som ska tilldelas ett makro.  
%PRODUCTNAME  
Om du väljer det här alternativet utförs det tilldelade makrot alltid när den valda händelsen uppträder, oberoende av dokumentet.  
Men detta gäller bara för globala makron.  
Makron som är bundna till dokument utförs bara när motsvarande dokument är laddat.  
Dokument  
Om du markerar alternativet Dokument utförs det tilldelade makrot bara vid en händelse, om det dokument som innehåller makrot är aktivt.  
Ett makro som du tilldelar händelsen Öppna dokument fungerar t.ex. som ett autostartmakro.  
Makron  
I området Makron visas i den vänstra listrutan de bibliotek och moduler som är tillgängliga och som innehåller dina makron.  
Om du klickar på plustecknet framför en post visas de underordnade posterna.  
Om du klickar på minustecknet döljs de underordnade posterna igen.  
De olika makrona är uppdelade i två områden som vart och ett är märkta med namnet på den översta posten i listrutan.  
I det andra finns globala makron som är dokumentoberoende.  
I den högra listrutan finns de makron som är tillgängliga för den modul som du valt i den vänstra listrutan.  
Tilldelningen sker enligt formatet "Subname(Bibliothekname.Modulname)".  
Programmeringsspråk  
I listrutan väljer du vilken typ av makron du vill integrera.  
Tilldela  
Den här kommandoknappen tilldelar makrot som är markerat i området Makron den händelse som är markerad under Händelse.  
Upphäv  
Rättstavning  
Här startar du rättstavningskontrollen med motsvarande kommando på undermenyn samt startar och stänger av den automatiska kontrollen.  
Kontrollera...  
Automatisk stavningskontroll  
Nytt fönster  
Med det här kommandot öppnar du ytterligare ett fönster för visning av den aktuella aktiviteten.  
När du har öppnat det nya fönstret visas det som ytterligare aktivitet.  
Innehållet i det nya fönstret visas först som en ny vy av det aktuella dokumentet.  
Ändringarna övertas alltid i dokumentets övriga fönster.  
Dokumentlista  
Detta gäller även för delade aktivitetsfönster.  
Det dokumentfönster som för närvarande visas markeras med en punkt framför namnet.  
Registrering  
Registreringen av %PRODUCTNAME sker online via vår registreringswebbsida.  
Registreringsdialogruta  
Andra gången du startar %PRODUCTNAME visas registreringsdialogrutan automatiskt med följande alternativ:  
Registrera nu öppnar vår registreringswebbsida i din standardwebbläsare.  
Registrera senare visar registreringsdialogrutan igen efter sju dagar.  
Om du väljer Registrera aldrig visas registreringsdialogrutan inte mer.  
Om du väljer Jag är redan registrerad visas registreringsdialogrutan aldrig mer.  
Använd det här alternativet om du t.ex. installerar om ditt %PRODUCTNAME efter registreringen.  
Du kan gå till registreringswebbsidan i din standardwebbläsare när du vill via Hjälp - Registrering.  
Lösenord  
I den här dialogrutan definierar du ett lösenord.  
Lösenord  
Ange ett lösenord som innehåller minst fem tecken i fältet Lösenord.  
Bekräfta  
Mata in samma lösenord en gång till för att bekräfta det.  
Upphäv lösenordsskydd  
När du öppnar dokumentet nästa gång måste du ange lösenordet.  
Om du anger fel lösenord går dokumentet inte att öppna.  
Inte ens våra programmerare kan då hjälpa dig.  
Definiera huvudlösenord  
I den här dialogrutan definierar du ett huvudlösenord för åtkomst till en lösenordsfil.  
En del lösenord kan sparas i %PRODUCTNAME.  
Beroende på sammanhanget kan du antingen spara ett lösenord så länge den aktuella %PRODUCTNAME -sessionen pågår eller så sparas det permanent i en fil.  
Lösenord för åtkomst till WebDAV-tjänster och FTP sparas permanent, om du markerar rutan Spara lösenord i motsvarande dialogrutor och tilldelar ett huvudlösenord.  
Om du inte tilldelar något huvudlösenord sparas bara lösenorden så länge den aktuella %PRODUCTNAME -sessionen pågår.  
Om du sparar permanent i en fil spärras filen med huvudlösenordet.  
Första gången du använder ett lösenord som har sparats permanent i en ny %PRODUCTNAME -session blir du automatiskt först ombedd att ange huvudlösenordet.  
Om du matar in det korrekt är alla lösenord som har sparats permanent kända i den aktuella %PRODUCTNAME -sessionen och du behöver inte ange dem igen.  
Huvudlösenord  
Ange ett huvudlösenord.  
Bekräfta huvudlösenord  
Ange samma huvudlösenord en gång till för att bekräfta det.  
Skriva ut fil direkt  
Om du klickar på ikonen Skriv ut fil direkt skrivs det aktiva dokumentet ut med de aktuella standardinställningarna.  
Dessa definierar du i dialogrutan Ställa in skrivare som du startar med menykommandot Skrivarinställning.  
Om du klickar på ikonen Skriv ut direkt när till exempel ett textområde eller ett grafikobjekt är markerat i ett öppet textdokument blir du tillfrågad om hela dokumentet eller enbart markeringen ska skrivas ut.  
Ritfunktioner  
Ikonen öppnar en utrullningslist med olika ritfunktioner.  
Information om att arbeta med ritfunktioner  
Ikon på utrullningslisten Ritfunktioner på verktygslisten:  
Visa ritfunktioner  
Urval  
Med den här ikonen markerar du ett objekt eller (med nedtryckt skifttangent) flera objekt, för att sedan flytta eller redigera dem gemensamt.  
Du kan också rita upp en urvalsram runt flera objekt.  
Samtliga objekt som ligger helt innanför urvalsramen markeras när du släpper musknappen.  
Om inte något ritobjekt är markerat och du väljer verktyget Urval, öppnas ritobjektlisten där du nu kan välja en förinställning för attributen för nya objekt.  
Välj en annan färg i stället för "Blå 7", t.ex. "Röd 7", och rita därefter flera rektanglar.  
De nya rektanglarnas standardfärg är "Röd 7"  
Linje  
Så här ritar Du en rak linje.  
Släpp musknappen.  
Om Du håller skifttangenten nedtryckt när Du drar infogas linjen bara i 45 graders vinkel.  
Om Du dubbelklickar på den färdiga linjen kan Du skriva in en text som orienterar sig efter linjen.  
Texten följer linjen i den riktning som Du har dragit den.  
Rektangel  
Med hjälp av denna ritar Du en rektangel, och med nedtryckt skifttangent ritar Du en kvadrat.  
Visa på den plats där kvadraten ska börja och dra musen med nedtryckt musknapp till motsatt hörnpunkt.  
Släpp musknappen.  
Du kan ändra rektangelns hörnrundning interaktivt, om du har aktiverat läget Redigera punkter.  
Ellips  
Med hjälp av denna ritar Du en ellips, och med nedtryckt skifttangent ritar Du en cirkel.  
Peka på den plats där ellipsen ska börja och dra musen med nedtryckt musknapp till motsatt slutpunkt.  
Släpp musknappen.  
Polygon  
Klicka här om du vill rita en polygon.  
Definiera de båda första punkterna genom att hålla ner musknappen och dra en linje.  
Klicka nu på varje ytterligare punkt i polygonen.  
Varje ny punkt förbinds automatiskt med föregående punkt.  
För att sluta polygonen dubbelklickar du på den första punkten.  
En linje dras från den sista punkten till den första och sluter polygonen.  
Om Du håller skifttangenten nedtryckt när Du ritar infogas de nya punkterna bara i 45 graders vinkel.  
Du kan ändra polygonens punkter interaktivt, om du har aktiverat läget Redigera punkter.  
Bézier  
Klicka på den här ikonen om du vill definiera en fri Beziérkurva.  
Nu kan du definiera en kurva i dokumentet genom att fastlägga tre punkter.  
Den första punkten är stället där du trycker ned musknappen.  
Håll ner musknappen och dra sedan till den andra punkten.  
Släpp musknappen.  
Klicka nu på den tredje punkten.  
När du klickar på den tredje punkten beräknar %PRODUCTNAME Bézierkurvan genom de tre punkterna och visar dem.  
Du avslutar kurvan genom att dubbelklicka.  
Om du håller ner Alternativ Alt -tangenten, avslutas kurvan också stängs kurvan.  
Frihand  
Så här ritar du en linje på frihand.  
Klicka där du vill att frihandslinjen ska börja och dra linjen som du vill ha med nedtryckt musknapp.  
När du släpper musknappen skapas linjens slutpunkt.  
Om du ritar ett slutet objekt, d.v.s. om du drar linjens slutpunkt till startpunkten, fylls ytan med den förvalda färgen.  
Cirkelbåge  
Klicka här om du vill rita ellipsbåge, håll ner skifttangenten om du vill rita en cirkelbåge.  
Sätt muspekaren i kanten av en tänkt ellips.  
Tryck på musknappen, håll ner den och rita upp ellipsen till önskad storlek.  
Släpp musknappen.  
Mellan centrum och ellipskonturen framträder nu en linje som följer varje musrörelse.  
Flytta centrumlinjen med musen till den önskade ellipsbågens start - eller slutpunkt och klicka.  
Centrumlinjen tas bort.  
Bestäm ellipsbågens storlek med musen och klicka.  
Ellipssektor  
Klicka här om du vill rita en ellipssektor, håll ner skifttangenten om du vill rita en cirkelsektor.  
Sätt muspekaren i kanten av en tänkt ellips.  
Tryck på musknappen, håll ner den och rita upp ellipsen till önskad storlek.  
Mellan centrum och ellipskonturen framträder nu en linje som följer varje musrörelse.  
Flytta centrumlinjen med musen till den önskade ellipssektorns start - eller slutpunkt och klicka.  
Centrumlinjen tas bort.  
Bestäm ellipssektorns storlek med musen och klicka.  
Cirkelsegment  
Klicka här om du vill rita ett ellipssegment, håll ner skifttangenten om du vill rita cirkelsegment.  
Sätt pekaren i kanten av en tänkt ellips.  
Tryck ner musknappen och rita med nedtryckt musknapp upp ellipsen till önskad storlek.  
Mellan centrum och ellipskonturen framträder nu en linje som följer varje musrörelse.  
Flytta centrumlinjen med musen till det önskade ellipssegmentets start - eller slutpunkt och klicka.  
Centrumlinjen tas bort.  
Bestäm ellipssegmentets storlek med musen och klicka.  
Text  
Klicka här om du vill definiera en textram där du kan skriva in text.  
Rita upp en rektangel genom att dra från det ena hörnet av rektangeln till det motsatta hörnet med nedtryckt musknapp.  
När du släpper musknappen visas begränsningen för textramen, som enligt standardinställningarna inte har någon synlig eller utskrivbar ram. (Men du kan ändra detta om du vill).  
Nu kan du börja skriva in text direkt.  
Den här texten kan du t.ex. rotera eller skala som grafikobjekt med hjälp av kommandona på formatmenyn.  
Klicka slutligen utanför inramningen om du vill återvända till den normala texten i dokumentet.  
Du kan ändra textramens hörnrundning interaktivt, om Du har aktiverat läget Redigera punkter.  
Animerad text  
Klicka på den här ikonen om du vill infoga animerad text i dokumentet.  
Håll ner musknappen och rita upp den ruta där den animerade texten ska röra sig.  
Med den här ikonen infogar du en animerad text i dokumentet.  
Håll ner musknappen och rita upp den ruta där den animerade texten ska röra sig.  
Släpp musknappen.  
Området där den animerade texten ska röra sig visas som en linje.  
Skriv nu texten som ska användas som animerad text.  
Klicka till slut på valfri plats utanför inramningen.  
Under Format - Text - Animerad text hittar du olika effekter som du kan tilldela den animerade texten.  
Du kan bara överföra en animerad text i HTML-exportformaten %PRODUCTNAME Writer, MS Internet Explorer och Netscape Navigator 4.0 till ett HTML-dokument.  
Förklaring  
Med den här ikonen definierar du en förklaring med markeringspil.  
Sätt muspekaren där markeringspilen ska infogas (dit den ska peka).  
Tryck på musknappen och håll ner den.  
Förklaringsrutan visas vid pekaren.  
Dra markeringspilen med nedtryckt musknapp till önskad position.  
Släpp musknappen.  
Dubbelklicka i den markerade förklaringsrutan eller på förklaringsrutans kant och skriv in texten.  
Klicka till slut på en valfri plats utanför inramningen. (Vilken effekten blir när du dubbelklickar beror på vad du har valt under Verktyg - Alternativ - Presentation - Allmänt, Tillåt snabbredigering och Bara textområde kan markeras.)  
Du kan ändra förklaringens hörnrundning interaktivt, om du har aktiverat läget Redigera punkter.  
Vertikal förklaring  
Här definierar du en vertikal förklaring med markeringspil  
Vertikal text  
Här definierar du en textram där du kan skriva en text vertikalt.  
Formulärfunktioner  
Med Formulär -ikonen öppnar du en utrullningslist med element och funktioner som du använder för att skapa ett interaktivt formulär.  
Det går bara att öppna utrullningslisten genom att klicka normalt på ikonen om inget kontrollfält har infogats i dokumentet ännu.  
Om det däremot finns ett kontrollfält i dokumentet, måste du hålla ned musknappen lite längre när du klickar på Formulär -ikonen för att utrullningslisten ska öppnas.  
Om du klickar snabbt aktiverar du alltid det senast infogade kontrollfältet som visas som aktivt element på ikonen.  
Ikon på verktygslisten:  
Formulär  
Formulärfunktionerna är tillgängliga i text-, HTML-, tabell-, presentations - eller teckningsdokument i %PRODUCTNAME.  
Formulärfunktioner är t.ex. textfält där användaren kan mata in text eller kommandoknappar, som startar en viss funktion när användaren klickar på dem.  
De här formulärelementen kallas kontrollfält i %PRODUCTNAME.  
Du kan göra ett utkast till ett formulär genom att i dokumentet infoga de olika kontrollfält som du behöver till formuläret och definiera deras egenskaper.  
Ett formulär kan även länkas till en databas.  
Till fälten överförs då de data som ska matas in i databasen eller som ska hämtas och visas från databasen.  
När du utformar en webbsida kan du skapa formulär som HTML-dokument.  
Sådana formulär kan användas till att låta användare skriva in data som sedan skickas via Internet.  
I HTML-dokument kan du använda alla funktioner när du skapar formulär, men du kan bara exportera de formuläregenskaper som stöds i den HTML-version som du använder.  
Du väljer HTML-version för export under Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet.  
Formulärfunktionerna i den aktuella versionen av %PRODUCTNAME stöds inte av versioner med lägre nummer än 5.0.  
Vid import och export av äldre dokumentversioner som innehåller kontrollfält görs ingen konvertering.  
Formuläregenskaperna försvinner vid såväl export som import.  
Om du vill infoga ett visst formulärobjekt i dokumentet, klickar du på motsvarande ikon på utrullningslisten.  
Muspekaren visar då med ett hårkors att du kan rita upp objektet i dokumentet.  
Om du vill skapa ett kvadratiskt kontrollfält, håller du ner skifttangenten medan du ritar.  
Om du i formuläret vill infoga fält från fältlistan i en tabell eller en sökning, kan du dra dem från den öppna tabellen eller sökningen till formuläret.  
Ett fältkommando infogas i textdokument om du enbart drar och släpper, om du samtidigt håller ner Kommando Ctrl och Skift skapas ett formulärfält.  
När du har infogat ett formulärelementet i dokumentet, kan du tilldela det önskade egenskaper.  
Markera kontrollfältet och klicka på ikonen Kontrollfältegenskaper eller välj kommandot Kontrollfält på kontrollfältets snabbmeny.  
En dialogruta öppnas där du kan definiera egenskaperna.  
Du kan kopiera kontrollfält från ett dokument till ett annat genom att dra och släppa dem eller använda Urklipp.  
Därvid utvärderar %PRODUCTNAME de tre egenskaperna "Databas", "Datakälla" och "Typ av datakälla "hos kontrollfältet, så att det hamnar på rätt ställe i måldokumentets logiska formulärstruktur.  
Ett kontrollfält som visar t ex ett innehåll i adressboken kommer att göra det även efter kopiering till måldokumentet.  
Kontrollfältet inordnas automatiskt i måldokumentet, antingen i den befintliga formulärstrukturen eller på så sätt att en struktur skapas.  
Följande kontrollfält finns:  
Kommandoknapp  
Med den här ikonen skapar du en kommandoknapp.  
Den kan du använda till att få ett kommando utfört vid en viss händelse, t.ex. då användaren klickar med musen.  
Kommandoknappar kan vara försedda med text och / eller grafik.  
Alternativfält  
Med den här ikonen skapar du ett alternativfält.  
Där kan användaren välja ett av flera alternativ.  
Alternativfält som hänger ihop funktionsmässigt får samma namn (Namn - Egenskap).  
De förses vanligen med en grupperingsram.  
Kryssruta  
Med den här ikonen skapar du en kryssruta.  
En kryssruta används till att sätta på eller stänga av en funktion.  
Etikettfält  
Med den här ikonen skapar du ett fält för visning av text.  
De här etiketterna eller etikettfälten är bara till visning av fördefinierad text.  
Inga inmatningar görs i de här fälten.  
Grupperingsram  
Med den här ikonen skapar du en ram där flera kontrollfält optiskt förs samman till en grupp eller ett område.  
Du kan t.ex. förse kryssrutor eller alternativfält med en grupperingsram för att visa att de hör ihop.  
Om du infogar en grupperingsram i dokumentet startar AutoPilot gruppelement, som hjälper dig att skapa en alternativgrupp.  
Info: om du ritar en grupperingsram kring befintliga kontrollfält och vill markera ett kontrollfält i efterhand måste du först välja kommandot Placering - Längst bak på grupperingsramens snabbmeny.  
Därefter kan du markera ett kontrollfält om du håller ner Kommando Ctrl -tangenten när du klickar på kontrollfältet.  
Grupperingsramen är enbart till för den optiska presentationen.  
Alternativfälten grupperas funktionellt när du namnger dem:  
Om du vill gruppera dem anger du samma namn under alla alternativfältens Namn -egenskap.  
Textfält  
Med den här ikonen skapar du ett textfält.  
Det är inmatningsfält där användaren kan skriva text.  
Textfält i formulär visar data eller tar emot nya.  
Listruta  
Med den här ikonen skapar du en listruta.  
Där kan användaren välja en post i en lista.  
AutoPiloten hjälper dig att skapa kontrollfältet.  
Kombinationsfält  
Med den här ikonen skapar du ett kombinationsfält.  
Det rör sig om en listruta som användaren kan öppna.  
Med egenskapen "Bara läsning" kan du bestämma om användaren ska kunna göra inmatningar i fältet eller inte.  
Användaren kan välja bland posterna på listan.  
Om formuläret är länkat till en databas och den kopplingen redan är aktiv, visas automatiskt AutoPilot - kombinationsfält när kombinationsfältet har infogats i dokumentet.  
Grafisk kommandoknapp  
Med den här ikonen skapar du en kommandoknapp som visas som ett grafikobjekt.  
Förutom den grafiska presentationen har den här kommandoknappen samma egenskaper som vanliga kommandoknappar.  
Grafiskt kontrollfält  
Med den här ikonen skapar du ett grafiskt kontrollfält.  
Det är enbart till för att hämta bilder från en databas.  
Om du dubbelklickar på ett sådant fält i formulärvyn öppnas dialogrutan Infoga grafik där du kan infoga bilden.  
Det finns dessutom en snabbmeny (inte i utkastläget) med kommandon för att infoga och radera grafik.  
I formuläret kan bilder från en databank visas och - om det grafiska kontrollfältet inte är skrivskyddat - nya grafikobjekt infogas i databasen.  
I så fall måste kontrollfältet hänvisa till ett databasfält av typen Bild.  
Ange därför datafältet i egenskaperna för kontrollfält under fliken Data.  
Filurval  
Med den här ikonen skapar du en kommandoknapp för filurval.  
Datumfält  
Med den här ikonen skapar du ett datumfält.  
Om du länkar formuläret till en databas, kan datumvärdena i formuläret hämtas från den databasen.  
Om du ger datumfältet egenskapen "Öppna", kan användaren öppna en kalender för val av datum nedanför datumfältet.  
Detta gäller även för ett datumfält i ett tabellkontrollfält.  
Användaren kan enkelt redigera datumfält med hjälp av piltangenterna.  
Beroende på markörens placering ökas eller minskas värdena stegvis för datum, månad eller år.  
Särskild information om datumfält.  
Tidsfält  
Med den här ikonen skapar du ett tidsfält.  
Om du länkar formuläret till en databas, kan tidsvärdena i formuläret hämtas från den databasen.  
Användaren kan enkelt redigera tidsfält med hjälp av piltangenterna.  
Beroende på markörens placering ökas eller minskas värdena stegvis för timme, minut eller sekund.  
Numeriskt fält  
Med den här ikonen skapar du ett numeriskt fält.  
Om du länkar formuläret till en databas, kan de numeriska värdena i formuläret hämtas från den databasen.  
Formaterat fält  
Med den här ikonen skapar du ett formaterat fält.  
Det är ett textfält för vilket du kan ange hur in - och utmatningen ska vara formaterad och vilka gränsvärden som gäller.  
Ett formaterat fält har särskilda kontrollfältsegenskaper (Format - Kontrollfält).  
Valutafält  
Med den här ikonen skapar du ett valutafält.  
Om du länkar formuläret till en databas, kan innehållet i valutafälten hämtas från den databasen.  
Maskerat fält  
Med den här ikonen skapar du ett maskerat fält.  
Ett maskerat fält består av en inmatnings - och en teckenmask.  
Inmatningsmasken styr vilka data användaren kan mata in och teckenmasken styr det maskerade fältets status när formuläret laddas.  
Maskerade fält fungerar inte i HTML-format.  
Tabellkontrollfält  
Med den här ikonen skapar du ett kontrollfält för en databastabell.  
Den hjälper dig att skapa kontrollfältet.  
Tabellkontrollfältet är en tabellarisk vy av ett databasformulär.  
Det är till för att ge en snabb överblick av data.  
Om du länkar formuläret till en databas kan du i tabellkontrollfältet se de data som finns i datakällan.  
Med det här kontrollfältet kan du arbeta på samma sätt som med inmatningsmasken i ett vanligt databasformulär: du kan mata in data, radera dem, ändra dem och så vidare.  
Särskild information om tabellkontrollfält.  
Urval  
Med den här ikonen aktiveras respektive inaktiveras muspekarens markeringsläge.  
I markeringsläget kan du markera kontrollfält i formuläret så att de t.ex. kan redigeras.  
Lägg till fält  
Automatiskt kontrollelementfokus  
Om du klickar på den här ikonen fokuseras det första formulärobjektet när du öppnar dokumentet.  
Om den här funktionen inte är aktiverad fokuseras texten när dokumentet öppnas.  
Ordningsföljden för aktivering som du har definierat gäller.  
Kommandon på snabbmenyn  
Ett kontrollfälts snabbmeny  
I ett kontrollfälts snabbmeny hittar Du bl a följande kommandon:  
Ersätt med  
Visar en undermeny där du kan välja en kontrollfälttyp, som ska ersätta det markerade kontrollfältet.  
När du väljer en kontrollfälttyp omvandlas det markerade kontrollfältet till det nya.  
Så många egenskaper som möjligt övertas.  
Textfält  
Det markerade kontrollfältet omvandlas till ett textfält.  
Kommandoknapp  
Det markerade kontrollfältet omvandlas till en kommandoknapp.  
Etikettfält  
Det markerade kontrollfältet omvandlas till ett etikettfält.  
Listruta  
Det markerade kontrollfältet omvandlas till en listruta.  
Kryssruta  
Det markerade kontrollfältet omvandlas till en kryssruta.  
Alternativfält  
Det markerade kontrollfältet omvandlas till ett alternativfält.  
Kombinationsfält  
Det markerade kontrollfältet omvandlas till ett kombinationsfält.  
Grafisk kommandoknapp  
Det markerade kontrollfältet omvandlas till en grafisk kommandoknapp.  
Filurval  
Det markerade kontrollfältet omvandlas till en kommandoknapp för filurval.  
Datumfält  
Det markerade kontrollfältet omvandlas till ett datumfält.  
Tidsfält  
Det markerade kontrollfältet omvandlas till ett tidsfält.  
Numeriskt fält  
Det markerade kontrollfältet omvandlas till ett numeriskt fält.  
Valutafält  
Det markerade kontrollfältet omvandlas till ett valutafält.  
Maskerat fält  
Det markerade kontrollfältet omvandlas till ett maskerat fält.  
Grafiskt kontrollfält  
Det markerade kontrollfältet omvandlas till ett grafiskt kontrollfält.  
Formaterat fält  
Det markerade kontrollfältet omvandlas till ett formaterat fält.  
Särskilda egenskaper för ett formaterat fält  
Formatering:  
Du kan ställa in den här egenskapen genom att i dialogrutan Egenskaper: Formaterat fält  
I textfältet för denna kommandoknapp visas ett exempel.  
Du kan inte redigera exemplet i textfältet, men Du kan radera det.  
Då visar det formaterade fältet sitt innehåll så som det står i databasen i den tabell som är kopplad till det formaterade fältet, utan att något ändras i formateringen.  
Om det formaterade fältet inte är kopplat till en databas, gäller en standardtalformatering.  
Om det formaterade fältet är kopplat till ett textfält i en databas, behandlas inmatningar i detta fält som text.  
Om det formaterade fältet är kopplat till ett fält i databasen som kan visas som tal, behandlas inmatningar som tal. (Datum och tid behandlas också internt som tal.)  
Min. värde och max. värde:  
Här anger Du minsta och högsta värde för det formaterade fältet.  
För formaterade fält som är kopplade till ett textfält, har dessa båda värden och det därefter beskrivna standardvärdet ingen betydelse.  
Gränsvärdena bestämmer utmatningen av existerande data (Exempel:  
Min. värde står på 5, det kopplade datafältet innehåller heltalsvärdet 3.  
Max. värde står på 10, och Du skriver in 20.  
Inskrivningen korrigeras och 10 skrivs i databasen).  
Om fälten för Min. värde och Max. värde inte fylls i, görs ingen begränsning.  
Standardvärde:  
Detta värde används som standard för nya dataposter.  
Om Du öppnar ett dokument som innehåller ett formaterat fält med %PRODUCTNAME version 5.1 (i den fanns den här fälttypen inte ännu), läses det formaterade fältet som ett textfält där.  
Om Du sparar dokumentet i 5.1-versionen, blir det formaterade fältet till ett textfält permanent.  
Särskilda tips för datumfält  
I datumfälten används för tvåsiffriga årtal det gränsvärde som du väljer för hela %PRODUCTNAME under Verktyg - Alternativ - %PRODUCTNAME - Allmänt.  
Om du skriver in ett tvåsiffrigt årtal, som inte ligger inom det inställda området, visas det med fyra siffror så att du kan kontrollera det.  
Om 1930 har definierats som gränsvärde, och du skriver 2034, så visas med andra ord 2034 och inte 34.  
Det inställda gränsvärdet sparas tillsammans med varje dokument.  
Om du sparar ett dokument med gränsvärdet 1930 ändrat och öppnar det i en äldre version av %PRODUCTNAME, visas en varning att okända data kan gå förlorade.  
I den äldre versionen av %PRODUCTNAME gäller bara det tidigare gränsvärdet 1930.  
Särskilda tips för tabellkontrollfält  
Du kan konfigurera ett tabellkontrollfält, om Du vill visa dataposterna på motsvarande sätt.  
Du kan alltså definiera datafält för datavisning eller dataregistrering på samma sätt som för ett vanligt databasformulär.  
Text-, datum-, tids - och valutafält, numeriskt fält, maskerat fält, markerings - och kombinationsfält.  
Vid kombinerade tids - och datumfält skapas två kolumner automatiskt.  
Under det totala antalet dataposter visas antalet markerade rader inom parentes, om några är markerade.  
Om du vill infoga kolumner i tabellkontrollfältet, klickar du i sidhuvudet och öppnar snabbmenyn.  
Här visas följande kommandon:  
Infoga kolumn  
Visar en undermeny där Du kan välja ett datafält, som ska övertas i tabellkontrollfältet.  
Ersätt med  
Öppnar en undermeny där du kan välja ett datafält som ska ersätta datafältet som är markerat i tabellkontrollfältet.  
Radera kolumn  
Raderar den markerade kolumnen.  
Kolumn...  
Öppnar den markerade kolumnens egenskapsdialogruta.  
Om Du klickar på en kolumn i utkastläge, öppnas också kolumnens speciella dialogruta Egenskaper.  
Kolumnegenskaperna motsvarar i huvudsak Kontrollfältegenskaperna.  
Dessutom har Du tillgång till egenskapen för kolumnbredd här.  
Dölj kolumn  
Döljer den markerade kolumnen.  
Egenskaperna behålls.  
Visa kolumner  
Öppnar en undermeny, där du kan välja de kolumner som ska visas igen.  
Om du bara vill visa en kolumn klickar du på kolumnens namn.  
Bara de 16 första dolda kolumnerna visas.  
Om det finns fler dolda kolumner, öppnar du med hjälp av kommandot Fler dialogrutan Visa kolumner.  
Fler...  
Öppnar dialogrutan Visa kolumner.  
I dialogrutan Visa kolumner markerar du de kolumner som ska visas.  
Håll ner Skift - eller Ctrl-tangenten om du vill markera flera poster.  
Alla  
Om du vill visa samtliga kolumner, klickar du på Alla.  
Konfigurera tabellkontrollfältet med dra-och-släpp:  
Visa datakällvyn och dra de önskade fälten med musen från datakällvyn till tabellkontrollfältets sidhuvud.  
Då skapas en förkonfigurerad kolumn.  
Om du håller ner tangentkombinationen Skift+Ctrl när du kopierar en tabellkolumn till tabellkontrollfältets kolumnhuvuden genom att dra och släppa, visas en undermeny.  
Välj här typ för kolumnen som ska infogas i tabellkontrollfältet.  
Kontrollfältegenskaper  
Med det här kommandot öppnar du en dialogruta där du redigerar egenskaperna för det markerade kontrollfältet.  
Du kan bara öppna dialogrutan om du befinner dig i utkastläget och ett kontrollfält är markerat.  
Om du matar in data i dialogrutan Egenskaper bör du observera att det går att göra inmatningar på flera rader i öppningsbara kombinationsfält.  
Detta gäller alla fält där ett SQL-uttryck kan anges samt för egenskaper hos text - eller etikettfält.  
Du kan öppna dessa fält och skriva text i den öppnade listan.  
Följande tangentkombinationer finns för detta:  
Tangenter  
Effekt  
Alt+Nedåtpil  
Öppnar kombinationsfältet.  
Alt+Uppåtpil  
Stänger kombinationsfältet.  
Skift+Retur  
Infogar ny rad.  
Uppåtpil  
Placerar markören på raden ovanför.  
Nedåtpil  
Placerar markören på raden nedanför.  
Retur  
Avslutar inmatningen i fältet och placerar markören i nästa fält.  
Precis som med vanliga kombinationsfält kan du öppna och stänga listan genom att klicka på pilknappen i fältets högerkant.  
Men inmatningen går att göra antingen i den öppna listan eller i textfältet ovanför.  
Ett undantag är de egenskaper som kräver visning i form av en lista, t.ex. egenskapen Listposter, som kan anges för kontrollfälten Listruta och Kombinationsfält.  
Här kan du bara redigera posterna när listan är öppen.  
Allmänt  
Under den här fliken definierar du allmänna egenskaper för ett kontrollfält i formuläret.  
Av det skälet är nedanstående egenskaper inte tillgängliga för alla kontrollfält.  
Vid HTML-export exporteras alltid tillhörande standardvärden och inte de aktuella värdena.  
Standardvärden fastställs alltefter typ av kontrollfält med egenskaperna Standardvärde (t ex för textfält), Standardstatus (för kryssrutor och alternativfält) och Standardmarkering (för listrutor).  
Aktiverad  
Om ett kontrollfält har egenskapen "Aktiverad" inställd på Ja, kan användaren av formuläret använda kontrollfältet.  
Kontrollfältet visas då gråtonat i formuläret.  
Antal rader  
Här anger du hur många rader som ska visas i den öppnade listan.  
Den här inställningen fungerar bara om alternativet Ja har valts under "Öppningsbar".  
För kombinationsfält med egenskapen Öppningsbar kan du ange här hur många rader som ska visas i den öppnade listan.  
För kontrollfält som inte kan öppnas är det fältets storlek och teckenstorleken som avgör hur många rader som får rum.  
Typ av kommandoknapp  
Här definierar du genom att välja typ vilken åtgärd som ska utföras när användaren klickar på kommandoknappen.  
För en kommandoknapp definierar du genom att välja typ vilken åtgärd som ska utföras när användaren klickar på kommandoknappen.  
När användaren klickar på knappen kan detta exempelvis leda till att data skickas eller till att värdena i andra kontrollfält återställs till standardvärdena. (Respektive standardvärde definieras i egenskaperna för kontrollfält.)  
Det finns följande alternativ och åtgärder:  
Typ  
Åtgärd  
Push  
När användaren klickar på kommandoknappen utförs ingen åtgärd.  
Reset  
När användaren klickar på kommandoknappen återställs inställningarna i andra kontrollfält till fördefinierade standardvärden (Standardstatus, Standardmarkering, Standardvärde).  
Användaren har därmed möjlighet att återkalla ändringar som har gjorts i ett formulär och återgå till standardinställningarna.  
Submit  
Om användaren klickar på kommandoknappen skickas data som har matats in i andra kontrollfält i det aktuella formuläret.  
Mottagaradressen anges under URL i Formuläregenskaper.  
URL  
Om användaren klickar på kommandoknappen aktiveras en URL.  
Adressen anger du under URL.  
Under Ram kan du ange målram.  
De nämnda kommandoknapparna används i HTML-dokument.  
För databasformulär spelar egenskapen Typ ingen roll.  
Öppningsbar  
Här kan du ange om kombinationsfältet ska kunna öppnas (Ja) eller inte (Nej).  
Kombinationsfält kan ha egenskapen "Öppningsbar".  
När användaren klickar på den öppnas listan med posterna.  
Under Antal rader kan du definiera hur många rader som ska visas på den öppnade listan.  
Kombinationsfält som infogas som kolumner i ett tabellkontrollfält är normalt alltid öppningsbara.  
Justering  
Här kan du definiera justeringsalternativet.  
Många kontrollfält har egenskapen Justering.  
Du kan välja om texten ska vara vänsterjusterad, högerjusterad eller centrerad.  
För etikettfält gäller justeringen fältrubriken, för textfält själva innehållet och för kolumner i ett tabellkontrollfält gäller den innehållet i tabellfälten (data).  
För kommandoknappar gäller justeringen justeringen av ett grafikobjekt som du kan visa tillsammans med en text eller i stället för en text.  
Fyll automatiskt  
Här kan du definiera om funktionen AutoComplete ska kunna användas på kombinationsfältet.  
Du kan definiera om funktionen AutoComplete ska kunna användas på ett kombinationsfält.  
Om du väljer "Ja", kommer den text som användaren skriver in att fyllas ut med den närmast följande post på listan vars inledande tecken stämmer med inmatningen.  
Etikettfält  
Här väljer Du från vilken källa etiketten till kontrollfältet ska hämtas.  
Texten i etikettfältet förs in överallt där annars namnet på det underliggande databasfältet måste stå - alltså t ex i filternavigatorn, i sökdialogrutan och som kolumnnamn i tabellvyn.  
För alternativfält (radioknappar) kan bara texten i gruppramen användas som etikettfält.  
Den texten gäller alltså för alla alternativfält i samma grupp.  
Om Du klickar på kommandoknappen... bredvid textfältet så visas dialogrutan Urval etikettfält.  
Här väljer du ett kontrollfält på listan över kontrollfält.  
Ta bort markeringen från fältet ingen tilldelning, eftersom annars inget kontrollfält tilldelas som etikettfält.  
Med det här fältet kan Du upphäva kopplingen till ett etikettfält.  
Bredd  
Här anger Du bredden (i millimeter) på kolumnen i tabellkontrollfält.  
För kolumnerna i ett tabellkontrollfält anger Du här kolumnbredden.  
Måttenheten är millimeter.  
Datapostmarkör  
Här väljer Du om den första kolumnen ska visas med kolumnrubrik, där t ex den aktuella dataposten anges med en liten pil.  
Datumformat  
Här anger Du önskat format för datumangivelse.  
För datumfält anger Du här formatet för hur datumet ska skrivas.  
Detta sker oavsett i vilken form användaren har gjort inmatningen.  
Rotationsknapp  
Med alternativet Ja blir kontrollfältet ett rotationsfält med pilknappar.  
Numeriska fält, valutafält, datum - och klockslagsfält kan infogas som rotationsfält i formuläret.  
Trefaldig status  
Den här egenskapen avgör om en kryssruta förutom värdena SANN och FALSK även ska kunna visa värdet NOLL från en ansluten databas.  
Den funktionen är tillgänglig enbart om databasen tillåter NOLL-värdet, dvs innehåller datafält som kan anta de tre tillstånden SANN, FALSK och NOLL.  
Den här egenskapen är definierad bara för databasformulär, inte för HTML-formulär.  
Skriv ut  
Om kontrollfältet ska synas vid utskrift av dokumentet, markerar Du den här egenskapen.  
Inmatningsmask  
Här definierar Du inmatningsmasken, vilket innebär att Du genom att ange en teckenkod bestämmer vilken typ av tecken som kan skrivas i kontrollfältet.  
För maskerade fält kan Du med en teckenkod begränsa vilka typer av tecken som kan skrivas i kontrollfältet.  
Inmatningsmaskens längd avgör antalet möjliga inmaningspositioner.  
Om användaren matar in ett tecken som inte motsvarar masken, kommer hela inmatningen att förkastas när fältet lämnas.  
Du kan använda följande tecken vid definition av en inmatningsmask:  
Tecken  
Innebörd  
L  
En textkonstant.  
Den här positionen kan inte redigeras.  
I fältet visas det tecken som finns i motsvarande position i teckenmasken.  
a  
Här kan tecknen a-ö skrivas in.  
Om en versal skrivs, förvandlas den automatiskt till gemen.  
A  
Här kan tecknen A-Ö skrivas in.  
Om en liten bokstav matas in omvandlas den automatiskt till en stor bokstav.  
c  
Här kan tecknen a-ö och 0-9 anges.  
Om en stor bokstav matas in omvandlas den automatiskt till en liten bokstav.  
C  
Här kan tecknen A-Ö och 0-9 skrivas in.  
Om en gemen skrivs, förvandlas den automatiskt till versal.  
N  
Bara tecknen 0-9 kan skrivas in.  
x  
Alla utskrivbara tecken kan skrivas in.  
X  
Alla utskrivbara tecken kan skrivas in.  
Om en gemen skrivs, förvandlas den automatiskt till versal.  
För teckenmasken ""__.__.2000" definierar du t.ex. inmatningsmasken "NNLNNLLLLL ", om du vill att användaren bara ska kunna mata in fyra siffror för att ange datum.  
Formatkontroll  
För kontrollfält som innehåller formaterat innehåll (datum, klockslag o.s.v.) finns funktionen formatkontroll.  
Om formatkontrollen är aktiverad (Ja), kan användaren bara skriva in de tecken som är tillåtna för formatet.  
För ett datumfält godtas t.ex. bara siffror och datumavgränsare, medan inmatning av bokstäver ignoreras.  
Ram  
Här anger du för en kommandoknapp av typen "URL" den målram där den laddade URL-sidan ska visas.  
För kommandoknappar som laddar en URL (URL-typ) när användaren klickar på dem, anger du som målram den ram där den laddade sidan ska visas.  
URL-adressen anger du under URL.  
Här kan du välja en post från den lista som öppnas och bestämma i vilken ram det följande dokumentet ska laddas.  
Det finns följande möjligheter:  
Post  
Betydelse  
_blank  
Det följande dokumentet visas i en ny, tom ram.  
_parent  
Det följande dokumentet visas i en parent, alltså en överordnad ram.  
Om det inte finns någon parent, visas dokumentet i samma ram.  
_self  
Det följande dokument visas i samma ram.  
_top  
Det följande dokumentet visas i ett toppfönster, d.v.s. i den högsta ramen i hierarkin.  
Om utgångsramen redan är ett toppfönster visas dokumentet i samma ram.  
Den här egenskapen är av intresse för HTML-formulär; för databasformulär har den ingen betydelse.  
Grafik  
En grafisk kommandoknapp har en Grafik -egenskap.  
Här anger Du sökväg och filnamn för den grafik som ska visas på knappen.  
Om Du väljer grafikfilen med kommandoknappen... överförs sökväg och filnamn automatiskt till textfältet.  
Hård radbrytning  
Här kan du tillåta en hård radbrytning för ett flerradigt fält.  
För flerradiga textfält kan du tillåta en hård radbrytning.  
Den egenskapen får bara effekt om du under Flerradig också har valt "Ja".  
Hjälptext  
Här kan du skriva en valfri hjälptext, som visas som Tips-hjälp för kontrollfältet.  
Tips-hjälpen visar texten i användarläge när muspekaren flyttas över kontrollfältet.  
För kommandoknappar av URL-typ visas hjälptexten i stället för den URL-adress som har angetts under URL.  
Hjälp-URL  
På så sätt kan den hjälp som hör till ett kontrollfält visas.  
Om kontrollfältet är markerat och användaren trycker på F1-tangenten, öppnas hjälpen för kontrollfältet.  
Bakgrundsfärg  
Här kan du välja kontrollfältets bakgrundsfärg.  
För de flesta typer av kontrollfält kan du definiera en bakgrundsfärg.  
Om du klickar på egenskapsfältet Bakgrundsfärg, öppnas en lista där du kan välja bland flera färger.  
Alternativet "Standard" övertar systeminställningen.  
Om den färg du vill ha inte finns på listan, klickar du på kommandoknappen... och kan sedan själv definiera en färg i dialogrutan Färg.  
Horisontal rullningslist  
Här definierar du om textfältet ska förses med en horisontell rullningslist (Ja) eller inte (Nej).  
Textfält kan förses med en vertikal och en horisontell bildrullningslist.  
Om textfältet ska ha en horisontell rullningslist, väljer du "Ja" för egenskapen Horisontal rullningslist.  
Intervall  
Här kan du ange en steglängd för rotationsfält.  
För numeriska fält och valutafält kan du ange en steglängd med egenskaper "Rotationsfält".  
Om användaren klickar på pilknapparna till rotationsfältet höjs eller minskas värdet med intervallvärdet.  
Listposter  
Här definierar du de listposter som ska visas i dokumentet.  
Öppna listan och skriv texten.  
För listrutor eller kombinationsfält definierar du här de listposter som ska visas i dokumentet.  
Öppna fältet Listposter och skriv texten.  
Se även informationen om inmatning och tangentbordsstyrning.  
Den förinställda listposten anges i kombinationsfältet Standardmarkering.  
De listposter som matas in här kan bara användas i formuläret om alternativet "Värdelista" är valt under fliken Data under Typ av listinnehåll.  
Om det inte är själva listposterna utan tilldelade värden - som inte syns i formuläret - som ska skrivas i databasen eller skickas till mottagaren av webbformuläret, så kan listposterna tilldelas andra värden med hjälp av en värdelista (med t.ex. värden i en databas).  
Den värdelistan definieras under fliken Data.  
Välj "Värdelista" under Typ av listinnehåll och ange under Listinnehåll de värden (t.ex. fältinnehållet i ett datafält) som ska tilldelas motsvarande synliga listposter i formuläret.  
För att tilldelningen ska bli korrekt är ordningsföljden i värdelistan avgörande.  
En listpost som anges på fliken Data under Listinnehåll motsvarar taggen <OPTION VALUE=...>.  
Max. datum  
Här anger Du ett datum för datumfältet som användaren inte ska kunna överskrida.  
För datumfält kan Du ange ett datum som användaren inte ska kunna överskrida; dvs om användaren försöker ange ett senare datum så godtas det inte.  
Max. textlängd  
Här anger Du hur många tecken som maximalt får skrivas in.  
För text - och kombinationsfält anger Du hur många tecken som maximalt för skrivas in.  
Om den här egenskapen är odefinierad, har standardinställningen värdet noll.  
Om kontrollfältet är bundet till en databas och textlängden ska hämtas från databasens fältdefinition, kan Du här inte ange någon textlängd.  
Inställningarna hämtas från databasen bara om kontrollfältsegenskapen inte har definierats (tillståndet "obestämt").  
Max. värde  
Här anger Du ett värde för kontrollfältet som användaren inte ska kunna överskrida.  
Det betyder att ett högre värde än så inte godtas.  
För numeriska fält och valutafält kan Du genom att definiera ett maxvärde se till att ingen användare kan ange ett högre värde.  
Max. tid  
Här anger Du för tidsfältet ett klockslag som användaren inte ska kunna överskrida.  
För tidsfält kan Du genom att definiera ett visst klockslag se till att ingen användare kan ange ett senare värde.  
Det betyder att ett senare värde än så inte godtas.  
Multimarkering  
Här anger Du om det ska vara tillåtet att markera flera poster i kontrollfältet.  
För listrutor kan Du ange om användaren ska kunna markera flera poster.  
Flerradig  
Med den här egenskapen anger Du om kontrollfältet ska kunna hantera radbrytning, så att texten kan visas på flera rader.  
I text - och etikettfält kan texten visas på flera rader.  
Radbrytning görs då antingen med returtangenten eller sker automatiskt vid kontrollfältets högerkant.  
Som standard hanteras inte radbrytning.  
Om Du vill att det ska vara möjligt, anger Du alltså den här egenskapen.  
Minimidatum  
Här kan du ange ett datum som användaren inte får underskrida.  
För datumfält kan du ange ett datum som användaren inte får underskrida.  
Om användaren försöker ange ett tidigare datum så godtas det alltså inte.  
Minimivärde  
Det betyder att ett mindre värde än så inte godtas.  
För numeriska fält och valutafält kan Du genom att definiera ett minvärde se till att ingen användare kan ange ett lägre värde.  
Minimitid  
Här anger Du för tidsfältet ett klockslag som användaren inte ska kunna underskrida.  
Det betyder att ett tidigare värde än så inte godtas.  
Antal decimaler  
Här definierar hur många decimaler som ska visas med värdet.  
För numeriska fält och valutafält kan du definiera hur många decimaler som ska visas med värdet.  
Namn  
Här anges namnet på kontrollfältet.  
Varje kontrollfält har egenskapen Namn, med vilken fältet entydigt kan identifieras.  
Namnet visas i Formulär Navigator och det används även när kontrollfältet anropas i ett makro.  
Som standard finns redan ett namn infört som identifierar kontrollfältet med beteckning och nummer.  
Du kan ändra namnet om Du vill.  
Om Du arbetar med makron måste Du tänka på att namnen på kontrollfälten måste vara entydiga.  
Namnet är inte bara till för att entydigt beteckna ett kontrollfält utan används även till att gruppera olika kontrollfält som hör ihop funktionellt.  
Kontrollfält med identiska namn utgör en gruppering.  
Grupperade element kan Du visa på bildskärmen med hjälp av grupperingsramar.  
Navigationslist  
Här kan Du ange om navigationslisten ska vara synligt in i tabellkontrollfältets nederkant (Ja) eller inte (Nej).  
Du kan efter behov visa eller dölja den.  
Bara läsa  
Här anger Du om kontrollfältet ska vara skrivskyddat (Ja) eller kunna redigeras av användaren (Nej).  
Om ett kontrollfält har egenskapen "Endast läsa" är det skrivskyddat och användaren kan inte redigera det.  
Den här egenskapen kan ges till alla kontrollfält där användaren normalt har möjlighet att skriva.  
När det gäller ett grafiskt kontrollfält, vars grafik hämtas från en databas, innebär den här egenskapen att användaren inte kan införa något nytt grafikobjekt i databasen.  
Ram  
Här anger Du om kontrollfältets ram ska vara transparent, platt eller ha 3D-utseende.  
För kontrollfält som är försedda med ram anger Du med egenskapen Ram hur ramen ska visas i formuläret.  
Du kan välja mellan Transparent, Platt eller 3D.  
Ordningsföljd  
Egenskapen Ordningsföljd definierar i vilken ordningsföljd kontrollfälten ska fokuseras när användaren trycker på tabbtangenten.  
Om det finns flera kontrollfält i ett formulär, flyttas alltså fokus till nästa kontrollfält i ordningen när tabbtangenten trycks ner.  
Den ordningsföljd i vilken detta sker kan du ange med ett index under Ordningsföljd.  
Index för det första kontrollfältet som ska fokuseras är 1.  
Egenskapen Ordningsföljd finns inte för Dolda kontrollfält.  
Inte heller grafiska kommandoknappar och grafiska kontrollfält går att välja med tabbtangenten.  
Varje nytt fält får ett index som ökas med 1 jämfört med föregående.  
Om Du ändrar indexet för ett kontrollfält, uppdateras automatiskt indexen för de övriga.  
Element som inte kan aktiveras (Tabbstopp = Nej) tilldelas ändå ett indexvärde.  
De kontrollfältet hoppas dock över när tabbtangenten trycks ned.  
Du kan också ange indexen för olika kontrollelement i dialogrutan Aktiveringsordningsföljd.  
Referensvärde  
Här anger Du ett referensvärde för webbformulär som ska användas när formuläret skickas till en server.  
För databasformulär skrivs det här värdet i det databasfält som har tillordnats kontrollfältet.  
Du kan tillordna alternativfält eller kryssrutor ett referensvärde.  
När ett webbformulär skickas till en server, vidarebefordras referensvärdet dit.  
För databasformulär skrivs det här värdet i det databasfält som har tillordnats kontrollfältet.  
Referensvärde för webbformulär  
Det kan vara praktiskt att använda referensvärden om Du skapar ett webbformulär och vill att information om tillståndet hos ett kontrollfält ska överföras till en server.  
Om kontrollfältet markeras av användaren, skickas motsvarande referensvärde till servern.  
Om Du inte anger något referensvärde och användaren har markerat kontrollfältet, överförs värdet "ON" när formuläret skickas.  
Om Du har en kryssruta för alternativet "man" och en för kvinna "kvinna "och Du för kryssrutan "kvinna" har referensvärdet 1 och för "man "referensvärdet 2, så överförs värdet 1 till servern om användaren markerar fältet "kvinna" och värdet 2 om fältet "man "markeras.  
Om de två rutorna är grupperade, överförs för hela grupperingen värdet "ON" om någon av rutorna har markerats.  
Vid grupperingar bör Du därför vara noga med att definiera referensvärden om informationen "ON" inte räcker till för att ange kontrollfältets tillstånd.  
Referensvärden för databasformulär  
Exempel:  
Om Du har en gruppering av de 3 alternativen "under arbete", "klar" och "återremitteras", med referensvärdena "ToDo", "OK "respektive "ÅR", införs referensvärdet i databasen när användaren har markerat respektive alternativ.  
Standardstatus  
Med den här egenskapen anger Du om ett visst alternativ eller en viss markering ska vara inställd som standard.  
När dokumentet laddas antas detta fördefinierade tillstånd.  
Kontrollfältets tillstånd definieras av en post som Du anger här när användaren klickar på en kommandoknapp av typen Återställ.  
För alternativfält som är grupperade definierar egenskapen Standardstatus det tillstånd hos gruppen som ska motsvara standardinställningen.  
Standardmarkering  
Här definierar du vilken av listposterna som ska vara förvald.  
För en listruta definierar du med den här egenskapen vilken av listposterna som ska vara förvald.  
Vid laddning av dokumentet antas denna definierade status.  
Den första listposten har nummer 0, nästa 1 och så vidare.  
När användaren klickar på en kommandoknapp av typen Återställ definieras listrutans tillstånd av den post som väljs här.  
Standardvärde  
Med standardvärdet anger Du vilken post som ska införas som standard i kontrollfältet.  
Det värdet införs när t ex ett formulär öppnas eller när nya dataposter ska matas in.  
När användaren klickar på en kommandoknapp av typen Återställ definieras kontrollfältets tillstånd av en post som Du anger här.  
Särskilt för datum - och tidsfält visas som standard aktuellt datum respektive aktuellt klockslag, om inget annat standardvärde har definierats.  
Standardknapp  
Med den här egenskapen definierar du att den här kommandoknappen ska utlösas när användaren trycker på returtangenten.  
I en dialogruta eller ett formulär med flera kommandoknappar utlöses en av dem när användaren trycker på returtangenten.  
Om användaren har öppnat dialogrutan eller formuläret, och inte har utfört någon annan åtgärd ännu, är kommandoknappen med den här egenskapen standardkommandoknapp.  
Den egenskapen bör aldrig tilldelas fler än en enda kommandoknapp i dokumentet.  
I webbsidesformulär träffar Du på den här egenskapen hos t ex sökmasker.  
Detta är inmatningsmasker som innehåller ett textfält och en kommandoknapp av typen Submit.  
Sökbegreppen skrivs i textfältet och sökningen startas genom att man klickar på kommandoknappen.  
Om nu kommandoknappen är definierad som standardkommandoknapp, kan användaren helt enkelt efter inmatning av sökbegreppet trycka på returtangenten för att starta sökningen.  
Placera symbol framför  
För valutafält anger Du här om valutasymbolen ska visas framför eller bakom talet.  
Som standard placeras den bakom.  
Tabbstopp  
Egenskapen Tabbstopp anger om ett kontrollfält i ett formulär kan markeras med tabbtangenten.  
Följande alternativ finns:  
Standard  
Det här kontrollfältet beter sig så som man kan förvänta sig.  
Exempelvis markeras inte ett etikettfält som standard, däremot ett textfält.  
Nej  
När tabbtangenten trycks ned, hoppas kontrollfältet över och nästa i ordningen aktiveras.  
Det värde som har angetts under Ordningsföljd bibehålls.  
Ja  
Kontrollfältet kan markeras med tabbtangenten.  
Tusentalsavskiljare  
Om tusentalsavgränsare ska infogas automatiskt, väljer Du här alternativet Ja.  
För numeriska fält och valutafält anger Du här om tusentalsavgränsare ska användas.  
Rubrik  
Egenskapen Rubrik bestämmer kontrollfältets etikett och visas i formuläret.  
Om kontrollfältet har egenskapen Rubrik avgör den kontrollfältets etikett som visas i formuläret.  
För kolumner i ett tabellkontrollfält anger Du spaltrubrik respektive synlig beteckning på datafältet.  
Om Du skapar ett nytt kontrollfält, används som standard den fördefinierade beteckningen i egenskapen Namn som etikett på kontrollfältet.  
Därvid sätts beteckningen samman av kontrollfältnamnet och ett heltal som anger kontrollfältets nummer, alltså t ex CommandButton1.  
Med egenskapen Rubrik kan Du ge kontrollfältet en annan beteckning, så att etiketten beskriver fältets funktion.  
Ändra alltså den posten om Du vill ge kontrollfältet en meningsfull och för användaren synlig beteckning.  
Om du vill ha en rubrik på flera rader, öppnar du fältet med hjälp av pilknappen.  
Du kan nu mata in en radbrytning med tangentkombinationen Kommando +Ctrl +Retur.  
Egenskapen Rubrik fungerar enbart som etikett för ett formulärelement på den yta som är synlig för användaren.  
Om Du arbetar med makron bör Du observera att ett kontrollfält som ska köras alltid ska anropas med egenskapen Namn.  
URL  
Här anger Du för en kommandoknapp av typen "URL" den URL-adress som ska laddas när man klickar på knappen.  
För kommandoknappar av URL-typ anger Du under URL den webbadress som ska laddas när man klickar på knappen.  
Det kan gälla vilken måladress som helst: en fil, ett nytt formulär eller en webbplats på Internet.  
Om muspekaren i användarläge pekar på kommandoknappen, visas URL-adressen som Tips-hjälp om Du inte har angett någon annan hjälptext.  
Vertikal rullningslist  
Här anger Du om textfältet ska förses med en vertikal rullningslist (Ja) eller inte (Nej).  
Textfält kan förses med en horisontell och en vertikal rullningslist.  
Om det ska ha en vertikal rullningslist, väljer Du för egenskapen Vertikal rullningslist alternativet Ja.  
Valutasymbol  
Här anger Du ett tecken eller en teckenföljd för valutasymbolen.  
För valutafält kan Du ange valutasymbolen genom att med egenskapen Valutasymbol ange önskat tecken eller teckenföljd.  
Värde  
Här anger Du de data som ska överföras från dolda kontrollfält.  
För ett dolt kontrollfält kan Du under Värde ange de data som ska överföras från det dolda kontrollfältet.  
De data överförs tillsammans med formuläret när det skickas.  
Tecken för lösenord  
Om textfältet är avsett för inmatning av lösenord, anger du här ASCII-koden för det tecken som ska visas i stället för de tecken som användaren skriver in.  
När en användare skriver ett lösenord i ett textfält kan du bestämma vilket tecken som ska visas i stället för de tecknen som användaren skriver.  
Ange ASCII-koden för det önskade tecknet vid Tecken för lösenord.  
255.  
Vilket tecken som har vilken ASCII-kod kan Du se i dialogrutan för specialtecken (Infoga - Specialtecken...).  
Teckenmask  
Här definieras teckenmasken.  
Den är alltså alltid synlig när formuläret har laddats.  
Om ett fält är maskerat måste Du definiera en teckenmask.  
Den innehåller startvärdena och är alltid synlig när formuläret har laddats.  
Med hjälp av teckenkoden i inmatningsmasken bestämmer Du vilken typ av inmatning som användaren kan göra i det maskerade fältet.  
Teckenmaskens längd måste alltid vara lika med inmatningsmaskens längd.  
I annat fall kommer inmatningsmasken antingen att kapas eller fyllas ut med blanksteg till inmatningsmaskens längd.  
Teckenuppsättning  
Här kan du välja vilken teckenuppsättning som ska användas vid formatering av text i kontrollfältet.  
För kontrollfält som ska ta emot synlig text i formuläret eller som har en rubrik, kan du välja en teckenuppsättning som ska användas vid visning av texten i formuläret.  
Klicka då på kommandoknappen... så kan du ange teckensnitt i dialogrutan Teckensnitt.  
Den valda teckenuppsättningen används sedan för beskrivning av kontrollfält eller bestämmer hur inmatningarna ska visas i inmatningsfälten - eller listrutorna.  
När det gäller tabellkontrollfält avgör teckenuppsättningen hur data ska visas.  
Förutom teckensnittet kan du i dialogrutan Teckensnitt även ange färgen på texten i kontrollfältet.  
Radhöjd  
Här anger Du radhöjden i ett tabellkontrollfält i millimeter.  
Måttenheten är millimeter.  
Tidsformat  
Här anger Du önskat format för angivelse av klockslag.  
För tidsfält anger Du här formatet för hur klockslaget ska skrivas.  
Tilläggsinformation  
Här anger Du ytterligare information eller upplysande text om kontrollfältet.  
För varje kontrollfält kan Du här ange ytterligare information eller upplysande text.  
Programmeraren kan använda det här fältet till att lagra kompletterande information som ska användas i en programkod.  
Exempelvis kan det här fältet användas för utvärdering av variabler eller andra parametrar.  
Data  
Under den här fliken kan du tilldela det markerade formulärelementet en datakälla.  
För formulär med databaskoppling definieras den tillhörande databasen i Formuläregenskaper.  
Funktionerna för detta hittar du där under fliken Data.  
Inställningsmöjligheterna på fliken Data för ett kontrollfält är beroende av kontrollfältet i fråga.  
Du ser bara de alternativ som på ett meningsfullt sätt kan definieras för kontrollfältet.  
På fliken finns följande fält:  
Datafält  
Här anger Du det fält i formulärtabellen som kontrollfältets datainnehåll ska vara länkat till.  
För databasformulär kan Du länka enskilda kontrollfält till datafält i en databas.  
Det finns följande möjligheter:  
Fall 1:  
Det finns bara en tabell för formuläret.  
Under Datafält anger Du det fält i formulärtabellen vars innehåll ska visas.  
Fall 2:  
Kontrollfältet hör till ett underformulär som skapas genom SQL-sökning.  
Under Datafält anges det fält från SQL-satsen vars innehåll ska visas.  
Fall 3 (bara för kombinationsfält):  
För kombinationsfält anger du under Datafält i vilket fält i den aktuella formulärtabellen värden ska lagras som användaren matar in eller väljer. (De värden som visas på kombinationsfältets lista bestäms med en SQL-sats som läggs in under Listinnehåll.)  
Fall 4 (bara för listrutor):  
Formulärtabellen innehåller inte de data som ska visas utan en tabell som är länkad till formulärtabellen via ett gemensamt datafält.  
Om data i en tabell som är länkad till den aktuella formulärtabellen ska visas i en listruta, anger du under Datafält det fält i formulärtabellen som listrutans datainnehåll är länkat till, respektive det databasfält som styr visningen av data i formuläret.  
Detta datafält anger kopplingen till den andra tabellen när båda tabellerna kan länkas via ett gemensamt datafält.  
Oftast rör det sig här om ett datafält där entydiga identifikationsnummer lagras. (Det datafält vars innehåll ska visas i formuläret anges via en SQL-sats under Listinnehåll.)  
Listrutor använder referenser.  
De kan realiseras antingen med hjälp av länkade tabeller via SQL-satser (fall 4) eller genom värdelistor:  
Referenser genom länkade tabeller (SQL-satser)  
Om en listruta ska visa data från en databastabell som via ett gemensamt datafält är länkad till den tabell som formuläret är baserat på, så visas under Datafält länkfältet i formulärtabellen.  
Länkningen sker via en SQL-Select, som för det valda alternativet "Sql" eller "Sql (Native) "anges i fältet Listinnehåll under Typ av listinnehåll.  
Om t.ex. kundnamn (som förvaltas i tabellerna "Kunder") ska visas i formuläret (tillhörande tabell "Beställning"), kan SQL-satsen lyda på följande sätt:  
SELECT Kundnamn, Kundnr FROM Kunder,  
där "Kundnamn" är datafältet i den länkade tabellen "Kunder "och "Kundnr" är det fält i tabellen "Kunder "som är länkat till det fält i formulärtabellen som anges under Datafält.  
Referenser via värdelistor  
De definierar referensvärden.  
På det sättet pekar kontrollfältet i formuläret inte direkt på ett innehåll i databasfältet utan på värden som tillordnas via värdelistan.  
Om Du arbetar med referensvärden på en värdelista ser Du i formulärets datafält inte det innehåll som Du har angett under Datafält, utan tillordnade värden:  
Om Du på fliken Data under Typ av listinnehåll har ställt in alternativet "Värdelista" och under Listinnehåll har tillordnat varje synlig listpost i formuläret (som Du ställer in på fliken Allmänt) referensvärden, kommer de referensvärdena att sättas lika med datainnehållet i de angivna datafälten.  
Om ett referensvärde motsvarar ett datafältinnehåll, visas de tillhörande listposterna i formuläret.  
Bundet fält  
Här anger Du med ett index vilket fält i en tabell eller en SQL-sökning som fältet som anges under Datafält är länkat med.  
Möjliga värden är 0, 1, 2, 3 osv.  
Denna egenskap, som står till förfogande för listrutor, avgör vilket datafält i en länkad tabell som ska visas i formuläret.  
Om en listrutat i formuläret ska visa innehållet i en tabell som är länkad till formulärtabellen, anger Du i fältet Typ av listinnehåll om visningen ska bestämmas med ett SQL-kommando eller om (den länkade) tabellen ska användas.  
Med egenskapen Bundet fält anger Du med hjälp av ett index det datafält som sökningen eller tabellen i listrutan är länkad till.  
Möjliga värden är 0, 1, 2, 3 osv.  
Egenskapen Bundet fält kan bara användas i formulär som är länkade till flera tabeller.  
Om bara en tabell ligger till grund för formuläret, anges under Datafält direkt vilket fält som ska visas i formuläret.  
Om listrutan däremot ska visa data från en databastabell som via ett gemensamt datafält är länkad till den aktuella tabellen, så bestäms det länkade datafältet av egenskapen Bundet fält.  
Om Du under Typ av listinnehåll har valt t ex alternativet "SQL", är det SQL-kommandot som bestämmer vilket index som ska anges.  
Exempel:  
Om ett SQL-kommando enligt formatet "SELECT fält1, fält2 FROM tabellnamn" är angivet under Listinnehåll så gäller:  
Bundet fält  
Länk  
0  
Databasfältet "fält1" är länkat till det fält som anges under Datafält.  
1  
Databasfältet "fält2" är länkat till det fält som anges under Datafält.  
Om Du under Typ av listinnehåll har valt alternativet "Tabell", är det tabellstrukturen som avgör vilket index som ska anges.  
Exempel:  
Om en databastabell har valts under Listinnehåll gäller:  
Bundet fält  
Länk  
0  
Kolumn nr 1 i tabellen är länkad till det fält som anges under Datafält.  
1  
Kolumn nr 2 i tabellen är länkad till det fält som anges under Datafält.  
2  
Kolumn nr 3 i tabellen är länkad till det fält som anges under Datafält.  
Typ av listinnehåll  
Här anger Du vilka data listan ska fyllas med.  
För listrutor och kombinationsfält anger Du med hjälp av listinnehållets typ vilka data listan ska fyllas med.  
Med alternativet "Värdelista" visas i kontrollfältet alla poster som Du har angett i fältet Listposter på fliken Allmänt.  
För databasformulär kan Du arbeta med referensvärden (se ovan).  
Om innehållet i kontrollfältet hämtas från en databas, kan Du ange typen av datakälla med de andra alternativen.  
Exempelvis kan Du här välja mellan tabeller och sökningar.  
Listinnehåll  
För databasformulär bestämmer Du här datakällan till formulärelementets listinnehåll.  
För dokument utan databaskoppling fungerar det här fältet så att det definierar en värdelista.  
För databasformulär bestämmer datakällan posterna i listrutor och kombinationsfält.  
Alltefter vilken typ som väljs - t.ex. tabell eller sökning - kan du under Listinnehåll välja mellan olika datakällor i den mån de objekten finns i din databas.  
Du kan här välja mellan alla databasobjekt av den typ som du har valt under Typ av listinnehåll.  
Om du har valt typen "Värdelista", kan du när det gäller databasformulär arbeta med referenser (se ovan).  
Om visningen av kontrollfältet regleras av ett SQL-kommando, införs SQL-satsen här.  
Exempel på SQL-sats:  
För listrutor har en SQL-sats exempelvis formen  
SELECT fält1, fält2 FROM tabell,  
där "tabell" är den tabell vars data visas i kontrollfältets lista (listtabell). "fält1 "är det datafält som bestämmer de poster som visas i formuläret; dess innehåll visas i listrutan. "fält2" är det fält i listtabellen som är länkat till formulärtabellen (värdetabellen) via det fält som anges under Datafält när Bundet fält = 1 har valts.  
För kombinationsfält har en SQL-sats exempelvis formen  
SELECT DISTINCT fält FROM tabell,  
där "fält1" är ett datafält i listtabellen vars innehåll visas i kombinationsfältets lista, dvs det datafält som bestämmer vilka poster som ska visas i formuläret.  
Värdelistor för HTML-dokument  
För HTML-formulär kan Du föra in en värdelista under Listinnehåll.  
Då väljer Du alternativet "Värdelista" under Typ av listinnehåll.  
De värden som Du här anger visas inte i formuläret utan är till för att tillordna de olika synliga posterna i formuläret värden som ska föras över vid exempelvis en dataöverföring.  
De inmatningar som har gjorts under Listinnehåll motsvarar HTML-taggen <OPTION VALUE=...>.  
Om det i den markerade positionen på värdelistan finns en (icke-tom) text (<OPTION VALUE=...>) överförs denna, annars överförs den text som visas i kontrollfältet (<OPTION>).  
Programmet tolkar den inmatningen som en tom sträng och tillordnar den till aktuell listpost.  
Följande tabell visar sambandet mellan HTML, JavaScript och %PRODUCTNAME -fältet Listinnehåll för en listruta med namnet "ListBox1".  
Här betecknar "Item" en listpost som visas i formuläret:  
HTML-tagg  
JavaScript  
Post på kontrollfältets värdelista (listinnehåll)  
Överförs...  
<OPTION>Item  
Inte möjlig  
""  
...den synliga listposten ("ListBox1=Item").  
<OPTION VALUE=" värde ">Item  
ListBox1.options[ 0].value="värde "  
"värde"  
...det värde som har tillordnats listposten ("ListBox1=värde").  
<OPTION VALUE=" ">Item  
ListBox1.options[ 0].value=" "  
"$$$empty$$$"  
...en tom sträng ("ListBox1=").  
Tom teckensträng är NOLL  
Här anger Du hur en tom teckenföljd vid inmatningen ska behandlas.  
I annat fall (Nej) behandlas teckenföljden som ett (tomt) värde.  
Filterförslag  
Medan du utarbetar ditt formulär kan du för varje textfält ange egenskapen "Filterförslag" under fliken Data i egenskapsdialogrutan för formuläret.  
I sådana fält kan du då vid en senare sökning i filterläge välja alla förekommande fältinnehåll i ett kombinationsfält.  
Då kan du också bekvämt välja fältinnehåll med hjälp av AutoComplete.  
Använd den därför sparsamt.  
Händelser  
Under den här fliken kan du länka vissa händelser, som kan inträffa för ett formulärkontrollfält, med ett makro.  
Makrot eller händelseproceduren sätts då igång så snart händelsen inträffar.  
Då öppnas en dialogruta där du kan välja makrot.  
Beroende på kontrollfält kan olika händelser inträffa.  
Under fliken Händelser finns därför bara de händelser som är möjliga för det markerade kontrollfältet.  
Följande händelser är definierade:  
Innan utförande  
Den här händelsen inträffar innan en åtgärd utlöses genom att användaren klickar på kontrollfältet.  
När du klickar på en submit-kommandoknapp, utlöser du visserligen åtgärden "skicka"; däremot startar själva processen att skicka först när händelsen "Vid utförande" inträffar.  
Med "Innan utförande" har du en möjlighet att stoppa verkställandet.  
Om den metod som är länkad till den här händelsen returnerar FALSE, utförs aldrig "Vid utförande".  
Vid utförande  
Den här händelsen inträffar när en åtgärd startas.  
Om du t.ex. har en kommandoknapp av typen submit i formuläret, utgör överföringsprocessen åtgärden.  
Modifierad  
Den här händelsen inträffar om kontrollfältet förlorar fokus och innehållet i kontrollfältet har ändrats sedan kontrollfältet fokuserades.  
Text modifierad  
Den här händelsen inträffar när text i ett inmatningsfält skrivs in eller ändras.  
Status ändrad  
Den här händelsen inträffar när kontrollfältets status ändras.  
För en kryssruta eller ett alternativfält är det när en ny post väljs.  
Vid fokusering  
Den här händelsen inträffar när ett kontrollfält fokuseras.  
Vid fokusförlust  
Den här händelsen inträffar när ett kontrollfält förlorar fokus.  
Efter tangenttryck  
Den här händelsen inträffar när användaren trycker på en valfri tangent medan kontrollfältet är fokuserat.  
Händelsen kan exempelvis vara länkad till ett makro som kontrollerar inmatningen.  
Efter tangenttryck  
Den här händelsen inträffar om användaren släpper en valfri tangent medan kontrollfältet är fokuserat.  
Mus inom  
Den här händelsen inträffar när muspekaren befinner sig inom kontrollfältet.  
Musrörelse vid tangenttryck  
Den här händelsen inträffar när musen flyttas medan en tangent hålls ner.  
Detta är exempelvis fallet när du drar och släpper om det är så att en tilläggstangent avgör dra-och-släppläget (förflyttning eller kopiering).  
Musrörelse  
Den här händelsen inträffar när musen flyttas över kontrollfältet.  
Musknapp nedtryckt  
Den här händelsen inträffar när musknappen trycks ner medan muspekaren är placerad på kontrollfältet.  
Musknapp uppsläppt  
Den här händelsen inträffar när musknappen släpps upp, medan muspekaren är placerad på kontrollfältet.  
Mus utanför  
Den här händelsen inträffar när muspekaren befinner sig utanför kontrollfältet.  
Formuläregenskaper  
I formuläregenskaperna definierar du bl.a. datakällan och händelserna för hela formuläret.  
Allmänt  
Under den här fliken definierar du allmänna egenskaper för formuläret.  
Med formulär menas ett elektroniskt formulärblad med olika kontrollelement.  
Om Du skapar ett formulär för en webbsida, kan användaren mata in data där som sedan skickas över Internet.  
Data i ett formulärs kontrollelement överförs till en URL-adress och kan där bearbetas vidare.  
Namn  
Med det namnet identifieras formuläret i Formulär Navigator.  
URL  
Ange här vilken URL-adress dit data i det formulär som användaren har fyllt i ska överföras.  
Ram  
I det här fältet anger Du den målram där det laddade URL-innehållet ska visas.  
Sändingstyp  
Välj här vilken metod som ska användas vid överföring av data i det formulär som användaren har fyllt i.  
Vid Get-metoden överförs data i varje kontrollelement som miljövariabel.  
Strängen utvärderas av ett program på mottagarens server.  
Det skickas sedan till den angivna URL-adressen.  
Kodning vid sändning  
Välj här typen av kodning för dataöverföringen.  
Dataöverföring av kontrollfältsinformation  
Vid sändning av ett formulär beaktas alla kontrollfält som är tillgängliga i %PRODUCTNAME.  
Kontrollfältets namn överförs alltid, likaså i förekommande fall det tillhörande värdet.  
Vilket värde som överförs beror på det aktuella kontrollfältet.  
För textfält överförs den post som visas; för listrutor de markerade posterna; för kryssrutor och alternativfält tillhörande referensvärden om fälten är markerade.  
Hur den här informationen överförs beror av den valda överföringsmetoden (Get eller Post) och kodningen (URL eller Multipart).  
Om t ex Get-metoden och URL-kodning används, skickas värdepar enligt formatet <namn>=<värde>.  
Utöver de kontrollfält som är kända inom HTML finns andra att tillgå i %PRODUCTNAME.  
Observera dock när det gäller fält med bestämda talformat att det inte är de värden som visas som överförs, utan motsvarande värden i fast definierade standardformat.  
Följande tabell visar hur data i %PRODUCTNAME -specifika kontrollfält överförs:  
Kontrollfält  
Värdepar  
Numeriskt fält, valutafält  
Ett decimaltecken anges alltid som punkt.  
Datumfält  
Datumformatet överförs som fast format (MM-DD-YYYY) oavsett användarens lokala inställningar.  
Tidsfält  
Tidsformatet överförs som fast format (HH:MM:SS) oavsett användarens lokala inställningar.  
Maskerat fält  
Värdet i ett maskerat fält överförs som textfält; dvs det som överförs är det värde som visas i formuläret.  
Tabellkontrollfält  
Från tabellkontrollfältet överförs alltid de enskilda kolumnerna.  
Det som skickas är kontrollfältets namn, namnet på kolumnen och kolumnens värde.  
Vid Get-metoden med URL-kodning genomförs överföringen exempelvis enligt formatet <tabellkontrollfältets namn>.<kolumnens namn>=<värde>, där värdet beror på kolumnen.  
Händelser  
Under den här fliken kan du tilldela ett makro vissa händelser som kan inträffa för ett formulär.  
Ett underordnat formulär reagerar även på de händelser som inträffar för det överordnade formuläret.  
Det kan då vara praktiskt att länka en händelse till ett makro om Du alltid måste reagera på ett visst sätt på en viss process i formuläret.  
Tillordna därefter händelsen i fråga makrot.  
Då öppnas en dialogruta där Du kan välja makro.  
Det innebär att Du kan använda Dina egna dialogrutor för att beskriva följande åtgärder:  
visa ett felmeddelande,  
bekräfta en radering (av dataposter),  
söka efter parametrar,  
och kontrollera inmatningar när en datapost sparas.  
På så sätt kan Du, när Du raderar en datapost, visa en kontrollfråga, som t ex "Vill Du verkligen radera kunden xyz?".  
Nedan beskrivs alla händelser som är definierade för ett formulär och som kan länkas till ett makro.  
Innan återställande  
Den här händelsen inträffar innan ett formulär återställs.  
Det länkade makrot kan t.ex. förhindra den här åtgärden genom att returnera FALSE.  
Ett formulär återställs när ett av följande villkor uppfylls:  
Användaren klickar på HTML-kommandoknappen som är definierad som Reset-kommandoknapp  
I ett formulär, som är bundet till en datakälla, skapas en ny, tom datapost när t.ex. kommandoknappen Nästa datapost används i den sista dataposten.  
Efter återställande  
Den här händelsen inträffar när ett formulär har återställts.  
Innan uppdatering  
Den här händelsen inträffar innan kontrollfältets innehåll som har ändrats av användaren skrivs i datakällan.  
Det länkade makrot kan t.ex. förhindra den här åtgärden genom att returnera FALSE.  
Efter uppdatering  
Den här händelsen inträffar när kontrollfältets innehåll som har ändrats av användaren har skrivits i datakällan.  
Före sändning  
Den här händelsen inträffar innan data i formuläret skickas.  
Vid laddning  
Den här händelsen inträffar direkt efter ett formulär har laddats.  
Före omladdning  
Den här händelsen inträffar innan formuläret laddas om.  
Datainnehållet har inte förnyats ännu.  
Vid omladdning  
Den här händelsen inträffar direkt efter en omladdning av ett formulär.  
Datainnehållet har redan förnyats.  
Före avladdning  
Den här händelsen inträffar innan ett formulär laddas av, d.v.s. skiljs från sin datakälla.  
Vid avladdning  
Den här händelsen inträffar direkt efter en avladdning av ett formulär, d.v.s. när ett formulär har skiljts från sin datakälla.  
Bekräfta radering  
Den här händelsen inträffar så snart raderingen av data utförs i formuläret.  
Det länkade makrot kan t.ex. efterfråga en bekräftelse i en dialogruta.  
Före datapoståtgärd  
Den här händelsen inträffar innan den aktuella dataposten ändras, t.ex. genom redigering, radering eller infogning.  
Det länkade makrot kan t.ex. efterfråga en bekräftelse i en dialogruta.  
Efter datapoståtgärd  
Den här händelsen inträffar direkt efter ändring av aktuell datapost, t.ex. genom redigering, radering eller infogning.  
Före datapostväxling  
Den här händelsen inträffar innan den aktuella datapostvisaren ändras, t.ex. genom kommandoknappen Nästa datapost.  
Det länkade makrot kan t.ex. förhindra den här åtgärden genom att returnera FALSE.  
Efter datapostväxling  
Den här händelsen inträffar direkt efter ändring av aktuell datapostvisare, t.ex. genom kommandoknappen Nästa datapost.  
Fyll parametrar  
Den här händelsen inträffar när det finns parametrar, som måste fyllas i, i formuläret som ska laddas.  
Formulärets datakälla kan t.ex. vara följande SQL-kommando:  
SELECT * FROM address WHERE name=:name  
Här är :name en parameter som måste fyllas vid laddning.  
Parametern fylls automatiskt från ett överordnat formulär under förutsättning att det är möjligt.  
Om parametern inte kan fyllas, startas den här händelsen och ett länkat makro kan fylla parametern.  
Fel har uppstått  
Den här händelsen inträffar när ett fel inträffar vid åtkomst till datakällan.  
Händelsen är definierad för formulär, listrutor och kombinationsfält.  
Data  
Under den här fliken definierar du formuläregenskaperna för en databas som är kopplad till formuläret.  
Här kan du bestämma på vilken datakälla formuläret ska basera eller om dessa data får påverkas av den som använder formuläret.  
Förutom sorterings - och filterfunktioner hittar du här alla nödvändiga egenskaper, som behövs för att skapa ett underordnat formulär.  
Om formuläret baseras på en SQL-sats (se egenskap Datakälla), är filter - och sorteringsfunktionerna bara tillgängliga om SQL-satsen bara refererar till en tabell och det inte heller är skrivet i databasens Native-SQL.  
Databas  
Här definierar Du databasen som innehåller datakällan som formuläret ska referera till.  
Genom att klicka på kommandoknappen... öppnar Du dialogen Öppna där Du kan välja ut den önskade databasen.  
Datakälla  
Här bestämmer du vilken datakälla som ska användas för formuläret.  
Datakällan kan för det första vara en existerande tabell eller sökning, som redan skapats i databasen, för det andra kan den definieras genom en SQL-sats.  
Innan du anger en datakälla måste du först definiera den exakta typen i fältet Typ av datakälla.  
Formulär, som är tilldelade en databas och som Du skapat i databasens formulärbehållare med hjälp av kommandot Nytt - Formulär, tillhör alltid databasen.  
För dessa formulär kan Du inte ändra datakällan i efterhand.  
Det kan Du bara (och det behövs bara), om Du med hjälp av utrullningslisten Formulärfunktioner gör ett "normalt "dokument till ett formulär.  
Om du har valt alternativet "Tabell" eller "Sökning "under Typ av datakälla, visas alla befintliga datakällor av den valda typen i kombinationsfältet, det vill säga alla tabeller resp. sökningar som har skapats i den markerade databasen.  
Om du vill basera formuläret på en sökning, måste du först välja alternativet "Sökning" som typ av datakälla, för att du ska kunna ange en sökning som datakälla.  
I fältet Datakälla kan du även ange en SQL-sats, om du valt alternativet "SQL" under Typ av datakälla.  
Med hjälp av den här satsen kan du skapa en SQL-sökning som ska ligga till grund för formuläret, eller definiera ett underordnat formulär.  
Typ av datakälla  
Här väljer du om en redan befintlig databastabell eller -sökning ska utgöra datakälla eller om formuläret ska genereras utifrån en SQL-sats.  
Om du väljer "Tabell" eller "Sökning ", baseras formuläret på den tabell eller sökning som du anger under Datakälla.  
Om du vill skapa en ny sökning eller skapa ett underordnat formulär, måste du välja alternativet "SQL".  
Du kan skriva in satsen för SQL-sökningen eller det underordnade formuläret direkt i fältet Datakälla.  
Formuläret genereras då utifrån den angivna satsen.  
Analysera SQL-kommando  
Om du har valt SQL-kommando under datakälla, definierar du här om SQL-kommandot ska analyseras (ja) eller inte (nej).  
Filter  
Här kan Du ange önskat villkor för filtrering av data i formuläret.  
Filter anges enligt SQL-regler utan att WHERE-instruktioner används.  
Om Du exempelvis vill visa alla dataposter med förnamnet "Klas" i en adressbokstabell skriver Du:  
Förnamn = 'Klas' (varvid "Förnamn "är namnet på datafältet).  
Man kan också kombinera flera villkor:  
Förnamn = 'Klas' ELLER Förnamn 'Mikael 'visar alla dataposter med förnamnen Klas och Mikael.  
Filterfunktionen är tillgänglig i användarläget genom ikonerna AutoFilter och Standardfilter på formulärlisten.  
Sortering  
Här kan Du ange önskat villkor för sortering av data i formuläret.  
Sorteringsvillkor anges enligt SQL-regler utan att ORDER BY-instruktionen används.  
Om Du exempelvis vill sortera alla dataposter i en adressdatabas stigande efter förnamn och inom förnamnen en gång till efter efternamn, anger Du:  
Förnamn ASC, Efternamn DESC (om "Förnamn "och "Efternamn" är namnen på databasfälten).  
Respektive ikoner på formulärlisten kan användas för sortering i användarläge:  
Sortera stigande, Sortera fallande, Sortera....  
Lägg endast till data  
Här definierar Du om formuläret bara ska tillåta att nya data läggs till (Ja) eller om det inte bara är begränsat till den här egenskapen (Nej).  
Användaren får bara lägga till data eftersom redan befintliga dataposter inte är synliga.  
Navigation  
Här anger Du om navigeringsfunktionerna på formulärlisten i formulärets nedre kant ska kunna användas (Ja) eller ej (Nej).  
Alternativet "Överordnat formulär" är till för underformulär.  
Om Du väljer detta alternativ för ett underformulär, kan Du navigera via dataposterna i huvudformuläret, om markören befinner sig i underformuläret.  
Då ett underformulär är kopplat till huvudformuläret genom en 1:1-relation, är det ingen vits att navigera inom ett underformulär.  
Navigationen utförs alltid på det överordnade formuläret.  
Cykel  
Här kan Du definiera hur navigationen ska ske inom formuläret med hjälp av tabbtangenten.  
Om Du samtidigt trycker ned skifttangenten navigerar Du i motsatt riktning.  
Om Du trycker på tabbtangenten när Du kommit till det sista (resp. det första) fältet i formuläret kan det få olika effekter.  
Du kan närmare definiera hur Du styr via tangentbordet med hjälp av följande alternativ:  
Alternativ  
Betydelse  
Standard  
Om det finns en databasanslutning i formuläret, går Du, om Du lämnar det sista fältet med hjälp av tabbtangenten, som standard till nästa / föregående datapost (se Alla dataposter).  
Utan databasanslutning går Du till nästa / föregående formulär (se Aktuell sida).  
Alla dataposter  
Detta alternativ är bara relevant för databasformulär.  
Med hjälp av det sker navigeringen över alla dataposter.  
När Du lämnar det sista fältet i ett formulär med hjälp av tabbtangenten byts den aktuella dataposten ut.  
Aktuell datapost  
Även detta alternativ är bara relevant för databasformulär.  
Med hjälp av det sker navigeringen bara inom en aktuell datapost.  
När Du lämnar det sista fältet i ett formulär med hjälp av tabbtangenten bevaras den aktuella dataposten.  
Aktuell sida  
När Du lämnar sista fältet i ett formulär hoppar Du till första fältet i nästa formulär.  
Det är standard för HTML-formulär, därför är detta alternativ särskilt relevant för HTML-formulär.  
Lägg till data  
Här definierar Du om data kan läggas till (Ja) eller inte (Nej).  
Ändra data  
Här definierar Du om data kan ändras (Ja) eller inte (Nej).  
Radera data  
Här definierar Du om data kan raderas (Ja) eller inte (Nej).  
Länka från  
Om Du skapar ett underformulär, anger Du här det överordnade formulärets datafält, vilket är ansvarigt för synkroniseringen mellan huvud - och underformulär.  
Om Du vill skriva in flera värden, trycker Du efter varje inmatningsrad på Kommando Ctrl +Retur.  
Det underordnade formuläret baseras på en SQL -sökning, närmare bestämt en parametersökning.  
Om du anger ett fältnamn i fältet Länka från, läses fältets data från huvudformuläret till en variabel, som du måste ange i fältet Länka till.  
Med hjälp av en lämplig SQL-sats jämförs den här variabeln med data i den tabell, som det underordnade formuläret refererar till.  
Genom detta tillvägagångssätt bestäms slutligen visningen i det underordnade formuläret.  
Här följer ett exempel.  
Den databastabell som ligger till grund för formuläret kan exempelvis vara en kunddatabas ("Kunder"), där Du ger varje kund ett entydigt nummer som beteckning, nämligen ett datafält kallat "Kund_ID ".  
Beställningarna från en kund organiserar Du i en annan databastabell.  
Nu vill Du också att beställningarna för varje kund som Du skriver in i formuläret ska visas.  
Då skapar Du underformuläret och skriver vid Länka från in datafältet från kunddatabasen, med hjälp av vilket kunden entydigt kan identifieras, det vill säga "Kund_ID" (utan citattecken).  
Vid Länka till skriver Du in namnet på en variabel, som ska ta med data i fältet Kund_ID, exempelvis "x".  
Underformuläret ska nu för varje kund resp. kundnummer (Kund_ID -> x) visa motsvarande data från beställningstabellen ("Beställningar").  
Det går naturligtvis bara om varje beställning entydigt är tilldelad en kund i beställningstabellen.  
Det kan också ske genom ett fält med namnet "Kund_ID", men för att vi inte ska förväxla det med fältet från huvudformuläret antar vi helt enkelt att det kallas "Kund_Nr".  
Nu behöver vi bara jämföra "Kund_Nr" i tabellen "Beställningar "med "Kund_ID" i tabellen "Kunder ", vilket kan uppnås genom variabeln x exempelvis med följande SQL-sats:  
SELECT * FROM Beställningar WHERE Kund_Nr =: x (om underformuläret ska visa samtliga data från beställningstabellen)  
eller:  
SELECT Artikel FROM Beställningar WHERE Kund_Nr =: x (om underformuläret från beställningstabellen bara ska visa data från fältet "Artikel")  
Du kan antingen ange SQL-satsen i fältet Datakälla eller skapa en motsvarande parametersökning, med vars hjälp du skapar ett underordnat formulär.  
Länka till  
Om du skapar ett underordnat formulär anger du här den variabel där möjliga värden från formulärets överordnade fält kan placeras.  
Om det underordnade formuläret bygger på en existerande sökning, anger du här den variabel som du har definierat i sökningen.  
Om du skapar det underordnade formuläret med hjälp av en SQL-sats, som skrivs in i fältet Datakälla, anger du här den variabel som du använder i satsen.  
Du kan välja fritt när du definierar variabelnamnet.  
Om du vill skriva in flera värden, trycker du på Kommando Ctrl +Retur efter varje inmatningsrad.  
Om du vid Länka från angett exempelvis databasfältet "Kund_ID" som överordnat fält, anger du vid Länka till namnet på den variabel, där värdena från databasfältet "Kund_ID "ska läsas in.  
Om du nu med hjälp av denna variabel anger en SQL-sats i fältet Datakälla, visas motsvarande värden i det underordnade formuläret.  
Vad är ett underordnat formulär?  
Formulär skapas utifrån en databastabell eller en databassökning.  
De kan också användas för redigering av befintliga data, vilka finns sparade i den databastabell eller -sökning som ligger till grund för formuläret.  
Om Du behöver ett formulär som inte bara har åtkomst till data i en tabell eller sökning, utan också ska visa data från ytterligare en tabell, kan Du skapa ett så kallat underformulär i Ditt formulär.  
Detta underformulär kan exempelvis bestå av ett textfält, som tar med data från en andra databastabell.  
Ett underordnat formulär är alltså ingenting annat än en "tilläggskomponent till ditt huvudformulär". "Huvudformuläret" betecknas som "överordnat formulär ".  
Alla andra data, som administreras i andra databastabeller, skapas som tilläggskomponenter i form av underordnade formulär.  
Underordnade formulär behövs alltså när du vill ha tillgång till mer än en tabell i ett formulär.  
För varje ytterligare tabell behöver du ett underordnat formulär.  
Som användare märker Du alltså inte att det är ett underformulär i sig.  
Du ser bara ett formulär, i vilket Du kan mata in Dina data eller där existerande data visas.  
Det är alltså möjligt att med hjälp av ett formulär med underformulär skapa en enkel inmatningsmask, som är helt anpassad till användarens behov, oberoende av hur dessa data organiseras i databasen.  
Ordningsföljd för aktivering  
I denna dialogruta kan Du ändra den ordningsföljd i vilken du går mellan kontrollfälten med tabbtangenten.  
Om formulärelement infogas i ett dokument bestämmer %PRODUCTNAME automatiskt i vilken ordningsföljd du går från ett kontrollfält till ett annat med tabbtangenten.  
Varje nytt kontrollfält tillfogas automatiskt i slutet av denna följd.  
I dialogrutan Aktiveringsordningsföljd kan Du påverka denna ordningsföljd och anpassa den till Dina individuella önskemål.  
Mata in det önskade värdet under Ordningsföljd i kontrollfältets egenskapsdialogruta.  
Kontrollelement  
Här listas samtliga kontrollfält som finns i det aktuella formuläret och som du kan välja med tabbtangenten.  
Välj ett kontrollfält genom att markera det och placera det i den önskade positionen i tabb-ordningsföljden.  
Index mindre  
Genom att klicka på denna kommandoknapp flyttar Du det markerade kontrollfältet ett steg upp i tabb-ordningsföljden.  
Index större  
Genom att klicka på denna kommandoknapp flyttar Du det markerade kontrollfältet ett steg ned i tabb-ordningsföljden.  
Auto sortering  
Klicka på denna knapp om Du vill sortera kontrollfälten automatisk inför fokuseringen med tabbtangenten.  
Den automatiska sorteringen beror på kontrollfältens position i dokumentet.  
Fälturval  
Klicka på den här ikonen om du vill öppna ett fönster där du kan välja ett databasfält som ska läggas till i formuläret.  
I fälturvalsfönstret listas alla databasfält i tabellen (eller sökningen), som du har angett som datakälla under Formuläregenskaper.  
Klicka på fältet med musen och dra det till dokumentet samtidigt som du håller ner musknappen.  
Det skapas då ett motsvarande fält i dokumentet med en länk till databasen.  
När Du stänger av utkastläget ser Du att %PRODUCTNAME lagt in ett etiketterat inmatningsfält för varje inmatat databasfält, i vilket användaren kan fylla i data.  
Designläge  
Med den här ikonen sätter du på eller stänger av utkastläget.  
I utkastläget kan du utforma formulärlayouten.  
Om det här läget inte är aktivt kan du inte bearbeta några formulärelement.  
Den här funktionen använder du för att snabbt växla mellan utkast - och användarläge.  
När du utformar ett formulär kan du växla läge om du t.ex. vill kontrollera formulärets utformning så långt.  
Var medveten om funktionen Öppna i utkastläge.  
Om denna funktion är aktiverad öppnas dokumentet alltid i utkastläge, oberoende av i vilket läge det har sparats.  
Om Du inte vill att användaren ska kunna öppna det färdiga formuläret i utkastläge stänger Du av denna funktion.  
Om formuläret är länkat till en databas visas formulärlisten vid dokumentfönstrets nedre kant när Du stänger av utkastläget.  
Länken till databasen anger Du i formuläregenskaperna.  
Formulär-Navigator  
Här visas samtliga formulär och de underordnade formulär som har skapats för det aktuella dokumentet, tillsammans med sina kontrollfält.  
Formulär-Navigator ger dig inte bara en nödvändig överblick när du arbetar med flera formulär, utan har också olika funktioner som du kan använda för att redigera ett formulär.  
I Formulär-Navigator visas en lista över alla (logiska) formulär, som har skapats i dokumentet, tillsammans med sina respektive kontrollfält.  
Om ett formulär innehåller kontrollfält indikeras detta av ett plustecken framför respektive post.  
Klicka på plustecknet så visas listan över formulärelement.  
Markera ett eller flera kontrollfält och dra det till ett annat formulär.  
Du kan även redigera beteckningen i Navigator genom att klicka på en post och ändra beteckningen.  
När Du väljer ett kontrollfält i Formulär-Navigator genom att klicka med musen markeras respektive element i dokumentet.  
På så sätt kan Du bekvämt navigera i dokumentet.  
Om Du anropar en markerad posts snabbmeny listas ett flertal funktioner i Navigator:  
Nytt  
Med detta kommando ställer Du funktioner till förfogande, som Du kan använda för att lägga till nya komponenter till formuläret.  
Dessa funktioner kan Du bara använda när ett formulär markerats i Navigator.  
Formulär  
Med detta kommando skapar Du ett nytt formulär.  
Om en formulärpost markerats skapas ett nytt underformulär till det markerade formuläret.  
Skapar ett dolt kontrollfält i det markerade formuläret.  
Kontrollfältet är inte synligt på bildskärmen och är därför dolt för användaren.  
Syftet med ett dolt kontrollfält är att du ska kunna ta emot de data som också överförs när ett formulär skickas iväg.  
Det innehåller ytterligare information eller förklarande text som du kan ange via kontrollfältets speciella egenskaper när du utformar formuläret.  
I vanliga fall kan du kopiera kontrollfält (tangentkombinationerna Kommando Ctrl +C för att kopiera och Kommando Ctrl +V för att klistra in).  
När det gäller dolda kontrollfält kan du naturligtvis inte göra på det här viset, eftersom de inte är synliga i dokumentvyn.  
Men du kan kopiera dolda kontrollfält i Formulär-Navigator med dra-och-släpp: dra det dolda kontrollfältet med musen och håll samtidigt ner tangenten Kommando Ctrl.  
Målet kan vara vilket formulär som helst, även det formulär där det dolda kontrollfältet redan finns.  
Genom att dra och släppa kan du kopiera kontrollfält i samma dokumentet och mellan olika dokument:  
Öppna ytterligare ett formulärdokument och dra det dolda kontrollfältet från Formulär-Navigator till måldokumentets Formulär-Navigator.  
Håll därefter musen stilla ett ögonblick så att kontrollfältet kan kopieras till urklippet.  
Dra sedan kontrollfältet till det andra dokumentet.  
Om du vill ha en kopia i samma dokument håller du ner Ctrl-tangenten när du drar.  
Radera  
Raderar den markerade posten.  
Med denna funktion kan Du radera såväl enskilda formulärkomponenter som hela formulär genom att klicka med musen.  
Ordningsföljd för aktivering  
När formuläret är markerat hämtas dialogrutan Aktiveringsordningsföljd, i vilken du definierar indexen för fokusering av kontrollelementen med tabbtangenten.  
Egenskaper  
Dialogrutan Egenskaper för den markerade posten visas.  
Om kontrollfältet markerats visas dialogrutan för kontrollfältsegenskaper.  
HTML-filter och formulär  
I HTML-dokument kan Du nu använda alla händelser som hör till kontrollelement och formulär.  
Tidigare fanns det många händelser (t ex Focus-händelserna) som inte ledde till någon åtgärd.  
Numera importeras och exporteras de som ONFOCUS, ONBLUR osv för JavaScript och som SDONFOCUS, SDONBLUR osv för %PRODUCTNAME Basic.  
En händelse som är registrerad som XListener::method exporteras som  
SDEvent-XListener-method = "/ * event-code * /"  
XListener - och metodkomponenterna i detta alternativ är skiftberoende (dvs skillnad görs mellan gemener och versaler)!  
Händelsehanteringen när det gäller Controls realiseras via %PRODUCTNAME API.  
Om Du tilldelar en Control en händelse, anmäls ett objekt som "Listener" för en viss händelse internt till Control-objektet.  
För att detta ska kunna ske måste det anmälda objektet ha ett visst gränssnitt, t ex XFocusListener Interface om det ska kunna reagera på fokus-händelser.  
När händelsen inträffar, anropar Control-objektet en viss metod i Listener-Interface, t ex focusGained, så snart Control-objektet erhåller fokus.  
Det internt anmälda objektet anropar då den JavaScript - eller %PRODUCTNAME -kod som har tilldelats händelsen.  
HMTL-filtret använder nu just dessa Listener-Interfaces och metodnamn för att kunna importera och exportera valfria händelser.  
I stället för att anmäla en fokus-händelse med  
<INPUT TYPE=text ONFOCUS=" / * code * / "  
kan Du även anmäla den med  
<INPUT TYPE=text SDEvent-XFocusListener-focusGained=" / * code * / "  
På detta sätt kan valfria händelser anmälas - även sådana som inte finns i listrutorna.  
För att fastställa skriptspråket för händelserna kan Du skriva följande rad i dokumenthuvudet:  
<META HTTP-EQUIV=" content-script-type "CONTENT="... ">  
För CONTENT kan Du använda bl a "text / x-StarBasic" för %PRODUCTNAME Basic eller ett "text / JavaScript "för JavaScript.  
Om Du inte anger någonting används JavaScript.  
Vid export bestäms standardskriptspråket av den första modul som hittas i makro-administrationen.  
För händelser kan alltså bara ett språk per dokument användas.  
AutoPilot för tabellelement  
Om du infogar ett tabellkontrollfält i ett dokument, startar AutoPilot för tabellelement automatiskt.  
Här kan du bestämma interaktivt vilken information som ska visas i tabellkontrollfältet.  
Du kan förhindra att autopiloterna startas automatiskt med ikonen AutoPilot på / av.  
AutoPilot för tabellelement / listruta / kombinationsfält - Data  
Här väljer du den datakälla och tabell som formulärfältet refererar till.  
När du infogar formulärfältet i ett dokument som som redan är kopplat till en datakälla visas inte den här sidan.  
Datakälla  
I det här fältet väljer du datakällan som innehåller tabellen som du vill använda.  
Tabell  
I det här fältet väljer du tabellen.  
AutoPilot för tabellelement - Fälturval  
Här väljer du vilka fält som ska visas i tabellkontrollfältet.  
Utvalda fält  
Här visas de datafält som används i formulärfältet.  
AutoPilot för kombinationsfält / listruta  
Om du infogar ett kombinationsfält eller en listruta i ett dokument, startar en AutoPilot automatiskt.  
I den här AutoPiloten bestämmer du interaktivt vilken information som visas.  
Du kan ställa av den automatiska starten av autopiloterna med ikonen AutoPilot på / av.  
Autopiloterna för kombinationsfält och listrutor skiljer sig i det sista steget.  
Det ligger i det här kontrollfältets natur:  
Listrutor  
I listrutor kan användaren välja en post bland flera på listan.  
Dessa poster är lagrade i en databastabell och kan inte redigeras i listrutan.  
Den databastabell som innehåller de listposter som visas i formuläret är normalt inte den tabell som formuläret baseras på.  
Listrutor i ett formulär arbetar därför med referenser på så sätt att referenser som hör till de visade listposterna finns i formulärtabellen (värdetabellen) och förs även in som sådana i värdetabellen när användaren väljer en post på listan och sparar den.  
Via referensvärden kan listrutor visa data från en tabell (listtabell) som är länkad till den aktuella formulärtabellen.  
Därför möjliggör AutoPilot för listruta länkningen av två tabeller i en databas, så att kontrollfältet kan visa en detaljlista från ett databasfält som finns i en annan tabell än den tabell som formuläret gäller.  
I den andra tabellen genomsöks det önskade fältet efter fältnamnet (ControlSource), och sedan fylls fälten i med motsvarande värden.  
Om fältnamnet inte kan hittas, förblir listan tom.  
För fältnamn med bundna kolumner införs den första spalten i den andra tabellen utan att någon bekräftelse krävs.  
Om exempelvis en artikeltabell innehåller numret på en leverantör, kan listrutan visa leverantörsnamnet från leverantörstabellen via länken "Leverantörsnummer".  
På sidan Fältlänk frågar autopiloten om alla inställningar som behövs för länken.  
Kombinationsfält  
I kombinationsfält kan användaren välja en post bland flera på listan eller själv skriva en text.  
De poster som finns på listan kan komma från valfri databastabell.  
De poster som användaren väljer eller anger för att de ska sparas kan sparas antingen i formuläret eller i en databas.  
Om de ska sparas i en databas, skrivs de in i den databastabell som formuläret är baserat på.  
Då får det inte finnas någon direkt koppling mellan den aktuella formulärtabellen och den tabell - listtabellen - vars värde ska visas i kombinationsfältet.  
I kombinationsfält används inte referenser.  
När användaren skriver in eller väljer ett värde och sparar det, införs detta värde i formulärtabellen.  
Eftersom det inte finns någon länk mellan formulär - och listtabellen, visas sidan Fältlänk inte här.  
Medan Du i en listruta kan välja bland poster på listan som är lagrade i listtabellen, kan Du i ett kombinationsfält dessutom skriva in egen text, som sparas i formulärets databastabell (värdetabellen) om Du så vill.  
Motsvarande alternativ finns inte för listrutor.  
Här kan Du ange om och var text som skrivs in i värdetabellen ska sparas.  
AutoPilot kombinationsfält / listruta:  
Tabellurval  
Här kan du bland de existerande tabellerna i databasen välja ut en tabell som innehåller det datafält vars innehåll ska visas som listposter.  
För listrutor anges här en tabell som kan länkas med den aktuella formulärtabellen.  
I så fall måste den länkade tabellen ha minst ett fält gemensamt med tabellen i det aktuella formuläret, så att det kan bildas en entydig relation.  
För kombinationsfält måste det inte finnas någon relation mellan formulärtabellen och den tabell som innehåller de data som ska visas i kombinationsfältet.  
Tabell för listinnehåll  
I detta fält väljer Du den tabell som innehåller det datafält vars innehåll ska visas i kontrollfältet.  
I kontrollfältsegenskaper na visas den här angivna tabellen som en del av en SQL-sats i fältet Listinnehåll.  
AutoPilot kombinationsfält / listruta:  
Fälturval  
Här väljer du från den tabell som angetts på den föregående sidan det datafält vars innehåll ska visas i kombinationsfältet eller listrutan.  
Existerande fält  
Här visas alla datafält i tabellen som du har valt i föregående steg i AutoPilot.  
Visningsfält  
Här anger du det fält vars data ska visas i kombinationsfältet eller listrutan.  
I kontrollfältsegenskaper na visas det här valda datafältet som en del av en SQL-sats i fältet Listinnehåll.  
AutoPilot listruta:  
Fältlänk  
Här anger du via vilka fält värde - och listtabellen är länkade.  
Listtabellen är den tabell vars data ska visas i listrutan.  
De båda tabellerna måste länkas via ett gemensamt datafält och denna länk anger du på den här sidan i AutoPilot.  
Fältnamnen måste inte nödvändigtvis överensstämma (det beror på hur fältnamnen i de två tabellerna har definierats), men båda fält måste ha samma fälttyp.  
Fält från värdetabellen  
Här anger Du det datafält i det aktuella formuläret som ska sättas i relation med ett fält i den länkade tabellen.  
Klicka på det önskade datafältet i den nedre listrutan.  
I kontrollfältsegenskaper na visas det här angivna fältet under Data -fliken som post under Datafält.  
Fält från listtabellen  
Här anger Du det datafält i den länkade tabellen som står i relation med det angivna fältet i värdetabellen.  
Klicka på datafältet i den nedre listrutan.  
I kontrollfältsegenskaper na visas det här angivna fältet under Data -fliken som del av en SQL-sats under Listinnehåll.  
AutoPilot för kombinationsfält:  
Databasfält  
För kombinationsfält kan du antingen spara ett fälts värde i ett databasfält eller bara använda det för visning i formuläret.  
Detta är lämpligt för HTML-formulär där de värden som användaren matar in eller markerar ska överföras till en server.  
Vill du spara värdet i ett databasfält?  
Det finns 2 alternativ för att svara på denna fråga:  
Ja, i följande databasfält  
Välj detta alternativ om det värde som användaren matat in eller markerat i kombinationsfältet ska sparas i ett databasfält.  
Du kan välja mellan samtliga fält ur den databastabell som det aktuella formuläret tilldelats.  
I kontrollfältsegenskaper na visas det här angivna fältet i data -registret som post under datafält.  
Listruta  
Här väljer Du det datafält i vilket kombinationsfältets värde ska sparas.  
Nej, jag vill bara använda värdet för visning  
Med detta alternativ sparas kombinationsfältets värde inte i databasen utan bara i formuläret.  
Öppna i redigeringsläge  
Om det här kommandot är aktiverat så öppnas formuläret i utkastläge när dokumentet öppnas.  
Du kan sedan redigera formuläret ytterligare, men du kan t.ex. inte klicka på några kommandoknappar i formuläret eller välja poster ur listrutorna.  
Upphäv kommandot när formuläret är färdigutvecklat, och sparar sedan formuläret ännu en gång.  
När formuläret öppnas nästa gång, kan alla interaktiva formulärelement användas.  
Ifall dokumentet är skrivskyddat så ignoreras detta kommando, dvs utkastläget aktiveras inte automatiskt vid dokumentets öppnande.  
Detta gäller t ex för databasformulären eftersom dessa som standard alltid är skrivskyddade.  
Autopilot på / av  
Med den här ikonen bestämmer du om AutoPilot ska startas automatiskt när ett nytt kontrollfält infogas.  
Den här inställningen gäller för alla dokument.  
AutoPiloter för infogning av en listruta eller ett kombinationsfält, ett tabellelement och för grupperingsramar.  
Visa raster  
Visa raster  
Fäst mot raster  
Om du klickar på den här ikonen blir rastret magnetiskt och objektet justeras alltid vid nästa rasterpunkt när det flyttas.  
Fäst mot raster  
Hjälplinjer vid förflyttning  
Hjälplinjer vid förflyttning  
Navigator  
Om du klickar på den här ikonen visar respektive döljer du Navigator.  
Du kan också starta Navigator med Redigera - Navigator Redigera - Navigator Redigera - Navigator Redigera - Navigator Redigera - Navigator.  
Navigator på / av  
Stylist  
Den används till att tilldela och administrera formatmallar.  
Du kan också starta Stylist med hjälp av Format - Stylist.  
Varje program i %PRODUCTNAME har en egen Stylist.  
Det finns alltså en särskild Stylist för textdokument textdokument, för tabelldokument tabelldokument och för presentationer / teckningsdokument presentationer / teckningsdokument presentationer / teckningsdokument.  
Stylist på / av  
Använd mall  
Med det här alternativet kan du tilldela det aktuella stycket eller de markerade styckena respektive ett markerat objekt en formatmall.  
Det finns fler mallar under Format - Stylist.  
Här ser du samma mallar som i mallistan i Stylist om du har valt mallgruppen Använda mallar i mallområdet.  
Använd mall  
Teckensnittsnamn  
Här väljer du teckensnittsnamnet från listan eller skriver namnet på ett teckensnitt direkt.  
Du kan mata in flera teckensnitt efter varandra med hjälp av semikolon.  
I så fall använder %PRODUCTNAME nästa teckensnitt när de föregående teckensnitten inte är tillgängliga.  
Ändringen gäller för den markerade texten eller ordet där markören står.  
Om ingen text är markerad gäller teckensnittsnamnet för texten som matas in därefter.  
De fem senast valda teckensnitten visas i övre delen av kombinationsfältet om du har markerat rutan Teckensnittshistorik under Verktyg - Alternativ - %PRODUCTNAME - Vy Så snart du stänger dokumentet återställs den vanliga alfabetiska uppräkningen av de installerade teckensnitten.  
Teckensnittsnamn  
Teckensnittsnamn  
I %PRODUCTNAME visas bara de existerande teckensnitten om en skrivare är installerad som standardskrivare i systemet.  
Du kan definiera en skrivare som standardskrivare med hjälp av programmet spadmin.  
Information om hur du installerar en skrivare som standardskrivare finns i dokumentationen till operativsystemet.  
Namnen på teckensnitten visas formaterade i respektive teckensnitt om du markerar rutan Förhandsvisning i teckensnittslistor under Verktyg - Alternativ - %PRODUCTNAME - Vy.  
Om det visas ett felmeddelande när du startar %PRODUCTNAME som talar om att vissa teckenuppsättningar inte går att hitta, kan du installera dem i efterhand med hjälp av setupprogrammet i reparationsläge, om det är fråga om ett %PRODUCTNAME -teckensnitt.  
Om du inte vill eller kan installera ett teckensnitt i efterhand kan du gå förbi felmeddelandet när du startar %PRODUCTNAME.  
Markera helt enkelt rutan Deaktivera meddelande.  
Teckenstorlek  
Här kan du välja mellan olika teckenstorlekar eller skriva in en teckenstorlek.  
Teckenstorlek  
Teckenstorlek  
Textriktning från vänster till höger  
Här kan du definiera den horisontella textriktningen.  
Textriktning från vänster till höger  
Textriktning uppifrån och ned  
Här kan du definiera den vertikala textriktningen.  
Textriktning uppifrån och ned  
Minska indrag  
Med den här funktionen minskar du det vänstra indraget i det aktuella stycket till föregående tabulatorposition.  
Genom att klicka på den här ikonen minskar du indraget av cellinnehållet i de markerade cellerna.  
Om du tidigare har ökat indraget för flera markerade stycken kan du minska indraget för dem med det här kommandot.  
Cellinnehållet flyttas med det värde som du har ställt in under Format - Cell... - Justering.  
Minska indrag  
Om du klickar på ikonen Minska indrag och samtidigt håller ner Kommandotangenten Ctrl-tangenten flyttas indraget för det markerade stycket med det standardtabbavstånd som är inställt under Verktyg - Alternativ - Textdokument - Allmänt.  
Öka indrag  
Med den här funktionen ökar du det vänstra indraget för det aktuella stycket till nästa tabulatorposition.  
Genom att klicka på den här ikonen ökar du indraget av cellinnehållet i de markerade cellerna.  
Om flera stycken är markerade ökas indraget för alla.  
Cellinnehållet flyttas med det värde som är inställt under Format - Cell... - Justering.  
Öka indrag  
Om du klickar på ikonen Öka indrag och samtidigt håller ner Kommandotangenten Ctrl-tangenten flyttas indraget för det markerade stycket med det standardtabbavstånd som är inställt under Verktyg - Alternativ - Textdokument - Allmänt.  
Exempel:  
Med ett standardtabbavstånd på 2 cm flyttas indragen för två stycken med hjälp av funktionen Öka indrag på följande sätt:  
Ursprungligt indrag  
Ökat indrag  
Indraget ökat med hjälp av Kommandotangenten Ctrl-tangenten med  
0,25 cm  
2 cm  
2,25 cm  
0,5 cm  
2 cm  
2,5 cm  
Teckenbakgrund  
Om du klickar länge på den här ikonen öppnas en utrullningslist där du kan tilldela en text en bakgrund i färg.  
Om du klickar kort tilldelar du markerad text den aktuella bakgrundsfärgen eller så aktiveras symbolen för färgöverstrykning (färgburk).  
Det finns två olika metoder.  
Om du klickar på ikonen och håller ner musknappen visas en utrullningslist där du kan välja bland förinställda bakgrundsfärger.  
När du har valt en färg får det ord som markören står i en bakgrund med den valda färgen.  
Den valda färgen visas på ikonen.  
Om du däremot klickar snabbt på ikonen ändrar muspekaren utseende och ser ut som en färgburk.  
Under den här symbolen visas ett grått, lodrätt streck som du använder för att markera ett textområde på samma sätt som med markören.  
Det här området tilldelas då automatiskt den bakgrundsfärg som du har valt på utrullningslisten Teckenbakgrund.  
Funktionen är aktiv så länge ikonen Teckenbakgrund är intryckt eller tills du trycker på Esc-tangenten.  
Om Du markerar Transparent på utrullningslisten Teckenbakgrund återställer Du bakgrundsfärgen.  
Teckenbakgrund  
Bakgrundsfärg Styckebakgrund  
Med den här ikonen visas en utrullningslist där du kan välja bland förinställda bakgrundsfärger.  
Om du vill tilldela enstaka celler i en tabell en bakgrundsfärg räcker det med att du ställer markören i motsvarande cell och klickar på önskad färg på utrullningslisten Bakgrundsfärg.  
Bakgrundsfärg  
Bakgrundsfärg)  
Styckebakgrund  
Växla objektlist  
Med den här ikonen växlar du mellan flera objektlister.  
Den här funktionen går bara att använda om flera olika objektlister är tillgängliga för redigering.  
Växla objektlist  
Öka styckeavstånd  
Genom att klicka på den här ikonen ökar du det övre styckeavståndet stegvis.  
Öka styckeavstånd  
Det finns mer information under Format - Stycke - Indrag och avstånd.  
Minska styckeavstånd  
Genom att klicka på den här ikonen minskar du det övre styckeavståndet stegvis.  
Minska styckeavstånd  
Det finns mer information under Format - Stycke... - Indrag och avstånd.  
Inramning  
Här ändrar du inramningen av ett tabellområde objekt.  
Det kan t.ex. gälla inramningen av en textram, ett grafiskt objekt eller en tabell.  
Ikonen på objektlisten visas bara när du har markerat ett grafikobjekt, en tabell, ett objekt eller en ram.  
Om du vill tilldela en enstaka cell en bestämd inramning räcker det om du placerar markören i den önskade cellen och klickar på en inramning på utrullningslisten Inramning.  
När du infogar ett grafikobjekt eller en tabell är dessa inramade.  
Därefter klickar du på ikonen som innebär "Ingen inramning" på utrullningslisten Inramning.  
Utrullningslisten Inramning  
Det finns mer information i hjälpen till Format - Stycke - Inramning.  
På ytterligare ett ställe finns information om hur du t.ex. utformar en texttabell med hjälp av inramningsikonen.  
Linjestil  
Med den här ikonen öppnar du utrullningslisten Linjestil där du kan ändra linjestilen för inramningen av ett objekt.  
Det kan t.ex. röra sig om inramningen av en ram, ett grafikobjekt eller en tabell.  
Ikonen på objektlisten visas bara om ett grafikobjekt, en tabell, ett diagramobjekt eller en ram markerats.  
Linjestil  
Det finns mer information under Format - Stycke - Inramning.  
Ramlinjefärg  
Med den här ikonen öppnar du utrullningslisten Inramningsfärg där du kan ändra linjefärgen i inramningen av ett objekt.  
Ikonen på objektlisten visas bara om ett grafikobjekt eller en ram har markerats.  
Ramlinjefärg  
Det finns mer information under Format - Stycke - Inramning.  
Byt förankring  
växlar du mellan en förankring vid cellen och vid sidan med ikonen Byt förankring. Var objektet är förankrat visas i dess snabbmeny. öppnar du en popupmeny med ikonen Byt förankring där du kan välja mellan olika förankringar.  
Ikonen visas bara på objektlisten när ett objekt, t.ex. ett grafikobjekt, ett kontrollfält eller en ram har markerats.  
Du kan förankra ett objekt vid sidan, vid ett stycke, vid ett tecken eller t o m som ett tecken.  
Om objektet omges av en ram kan det även förankras vid ramen.  
Du kan förankra ett objekt vid sidan, vid ett stycke, vid ett tecken eller t o m som ett tecken.  
Det finns mer information om olika förankringsalternativ i hjälpen till Format - Förankring.  
Linjeslutsstil  
Med ikonen Linjeslutsstil öppnar du utrullningslisten Linjeslut.  
Med hjälp av ikonerna där definierar du stil för den markerade linjens ändar.  
Den här ikonen visas bara på objektlisten när du har skapat en teckning med ritfunktionerna och markerat den.  
Det finns mer information i hjälpen till Format - Linje - Linjeslut.  
Linjeslutsstil  
Objekt-rotationsläge  
Om ikonen är aktiv (intryckt) kan du rotera det markerade objekt eller objekten med musen.  
Markera först ett objekt, klicka på ikonen på objektlisten och rotera sedan det markerade objektet genom att dra med musen.  
Den här ikonen visas bara på objektlisten när minst ett ritobjekt är markerat.  
Det finns mer information i hjälpen till menykommandot Format - Position och storlek... - Rotation.  
Objekt-rotationsläge  
Justera objekt Justera objekt Justering  
Med den här ikonen öppnar du utrullningslisten Justering.  
Nu kan du ändra justeringen av ritobjektet.  
Ikonen på objektlisten visas bara när ett ritobjekt är markerat.  
Det finns mer information finns i hjälpen till menykommandot Format - Justering.  
Justera objekt Justera objekt Justering  
En nivå nedåt NivÃ¥ lÃ¤gre  
Den här ikonen flyttar ned de markerade styckena i hierarkin.  
Ikonen visas bara när markören står i en punktuppställning eller numrering.  
Den visas på verktygslisten när du är i dispositionsvyn.  
En nivå nedåt Nivå lägre  
En nivå uppåt NivÃ¥ uppÃ¥t  
Den här ikonen flyttar upp de markerade styckena i hierarkin.  
Den visas bara när markören står i en punktuppställning eller numrering.  
Den visas på verktygslisten när dispositionsvyn är aktiv.  
En nivå uppåt Nivå upp  
Flytta uppåt UppÃ¥t  
Det aktuella stycket (eller alla markerade stycken) flyttas ett stycke uppåt.  
Inom en numrering anpassas numren till den nya positionen.  
Ett stycke flyttas maximalt till gränserna för den aktuella punktuppställningen eller numreringen eller det "normala" området upp till nästa punktuppställning eller numrering.  
Ikonen på numreringsobjektlisten visas bara när markören står i en punktuppställning eller numrering.  
Ikonen visas på verktygslisten när du är i dispositionsvyn.  
Du aktiverar den här funktionen genom att trycka på Kommando Ctrl +Uppåtpil.  
Flytta uppåt Uppåt  
Flytta nedåt NedÃ¥t  
Det aktuella stycket (eller alla markerade stycken) flyttas ett stycke nedåt.  
Inom en numrering anpassas numren till den nya positionen.  
Ett stycke flyttas maximalt till gränserna för den aktuella punktuppställningen eller numreringen eller det "normala" området ned till nästa punktuppställning eller numrering.  
Ikonen på numreringsobjektlisten visas bara när markören står i en punktuppställning eller numrering.  
Ikonen visas på verktygslisten när du är i dispositionsvyn.  
Du aktiverar den här funktionen genom att trycka på Kommando Ctrl +Nedåtpil.  
Flytta nedåt Nedåt  
Punktuppställning på / av  
Genom att klicka på den här ikonen förser du markerade stycken med punktuppställningstecken eller upphäver en punktuppställning.  
I dialogrutan Numrering / punktuppställning definierar du typ av punktuppställning.  
Du kan ändra strukturen med hjälp av ikonerna på numreringsobjektlisten.  
Du växlar till den här listen genom att klicka på pilknappen längst till höger på objektlisten.  
I Onlinelayout -läge är några av alternativen för numrering / punktuppställning inte tillgängliga.  
Avståndet mellan texten och den vänstra textramen kan Du ställa in i dialogrutan under Format - Stycke... genom att definiera vänsterindrag och förstaradsindrag.  
Du kan även lätt ställa in indragen med musen genom att dra i linjalen.  
Punktuppställning på / av  
Ladda URL  
I det här kombinationsfältet matar du in URL:en för dokumentet som du vill ladda.  
Du kan ange en ny URL eller välja en som redan har matats in. %PRODUCTNAME omvandlar automatiskt filsökvägar till URL-skrivsättet.  
Om du vill ladda ett nytt dokument som har en liknande URL som det aktuella dokumentet redigerar du URL-posten i kombinationsfältet och trycker på returtangenten. %PRODUCTNAME hjälper dig genom att känna igen liknande inmatningar och ge förslag så att du ofta bara behöver mata in delar av en URL.  
Ladda URL  
Du kan flytta inmatningsfokus direkt till fältet Ladda URL med tangentkombinationen Kommando Ctrl +Skift+O.  
Om funktionslisten är placerad lodrätt så visas i stället för det långa kombinationsfältet ikonen Ladda URL.  
Om du klickar på den här ikonen öppnas dialogrutan Öppna.  
Ladda URL  
Ladda på nytt  
Med det här kommandot ersätts det aktuella dokumentet med den senast sparade versionen.  
Eventuella ändringar som du har gjort sedan du senast sparade dokumentet går förlorade.  
Först görs dock en säkerhetskontroll.  
Redigera fil  
Om den här ikonen är intryckt (men inte dold) eller om du väljer det här kommandot kan du redigera det aktuella dokumentet eller databastabellen.  
Men den här funktionen sätter du på eller stänger av redigeringsläget.  
Redigera fil  
På titellisten visas om dokumentet som du har öppnat är skrivskyddat.  
Det betyder att du t.ex. har öppnat det från en cd-rom eller en nätverksenhet där du inte har några skrivrättigheter, eller att någon annan i nätverket redan har öppnat dokumentet.  
Klicka på ikonen Redigera fil på funktionslisten.  
Du tillfrågas om du vill redigera en kopia av dokumentet.  
Bekräfta frågan.  
Du kan redigera och spara kopian där du har skrivrättigheter.  
Redigera data  
Med den här ikonen sätter du på och stänger av redigeringsläget för den aktuella databastabellen.  
Redigera data  
Redigering av databaser i nätverk  
Om du vill göra ändringar i en databas som används gemensamt så måste du ha de nödvändiga skrivrättigheterna.  
Om du redigerar en extern databas sparas inte ändringarna som du gör av %PRODUCTNAME utan skickas direkt vidare till databasen.  
Spara aktuell datapost  
Genom att klicka på den här ikonen på Databaslisten sparar du den aktuella dataposten i databastabellen.  
Änderingar av innehållet i en datapost sparas automatiskt så fort du väljer en annan datapost.  
Använd den här ikonen om du vill spara ändringar, men inte vill välja någon annan datapost.  
Stoppa laddning  
Om du håller ner Kommando Ctrl samtidigt avbryts all laddning som pågår.  
Stoppa laddning  
Dokumentinformation  
I det här fältet får du information om det öppnade %PRODUCTNAME Basic-dokumentet.  
Namnet på dokumentet, biblioteket och modulen skiljs åt med en punkt.  
Position i dokumentet  
I det här fältet ser du vid vilken position i dokumentet markören står.  
Först anges radnumret och därefter kolumnnumret.  
URL-namn  
I det här kombinationsfältet kan du tilldela en Internet-URL eller en fil ett namn.  
Du kan även skriva en söktext som överförs till en sökmotor.  
Du kan använda följande syntax vid textsökning:  
Star+Office  
Hittar alla sidor som någonstans innehåller orden / orddelarna "Star" OCH "Office ".  
Star,Office  
Hittar alla sidor som innehåller "Star" ELLER "Office.  
Star Office  
Hittar alla sidor som innehåller den här texten.  
Sådana ordkombinationer överförs direkt till önskad sökmotor på Internet.  
I de flesta fall behandlar sökmotorerna ordkombinationen som en ELLER-förbindelse och söker alltså efter sidor som innehåller minst ett av orden.  
Vissa sökmotorer gör åtskillnad mellan versaler och gemener.  
Om Du är osäker är det bäst att skriva in alla bokstäver som gemener.  
Alla Internet - sökmotorer stöder dock inte alla logiska kombinationer.  
Använd endast något av de här tre alternativen för kombination av sökbegrepp när du startar en sökning.  
URL-namn  
Samlingsbox till webbadresser  
Här kan du antingen skriva en URL eller infoga en URL genom att dra och släppa den från ett dokument.  
Du kan redigera URL:en och infoga den på textmarkörens position i det aktuella dokumentet genom att klicka på Länk.  
Ikonen Länk går bara att aktivera om det finns text i fältet URL-namn.  
Samlingsbox till webbadresser  
Länk  
Genom att klicka på den här ikonen infogar du en hyperlänk till den aktuella URL:en i dokumentet.  
URL:en hämtas då från Samlingsbox till webbadresser, namnet från kombinationsfältet URL-namn.  
När Du klickar på ikonen får Du upp en meny, där Du kan definiera om hyperlänken ska infogas som text eller knapp.  
Visa på ikonen Länk, tryck på musknappen och håll den nedtryckt ett ögonblick.  
En urvalsmeny visas, där Du kan välja mellan alternativen Som text eller Som knapp.  
Flytta pekaren till önskat alternativ och släpp musknappen.  
Hyperlänken visas då, beroende på vad Du har valt, antingen som text i färg och understruken eller som knapp.  
Länk  
Sök  
Genom att klicka på den här ikonen öppnar du en lista där du kan välja en av de definierade Internet-sökmotorerna.  
Sökordet hämtas från från kombinationsfältet URL-namn.  
Texten som ska sökas måste finnas i kombinationsfältet.  
Klicka på ikonen Sök och håll ner musknappen.  
Då öppnas en undermeny där du kan välja en sökmotor.  
Sökmotorer definierar du via Verktyg - Alternativ - Internet - Sökning.  
Sök  
Sökmotorlista  
Om du har valt en av sökmotorerna överför %PRODUCTNAME sökförfrågan till din webbläsare som sedan skapar Internetförbindelsen till sökmotorn och visar resultatet.  
Se även URL-namn.  
Ram  
Med den här ikonen väljer du målram (target frame) för den angivna URL:en.  
Om du klickar på den här ikonen öppnas en undermeny med de fördefinierade ramarna.  
Ram  
Hyperlänkdialogruta  
Med den här ikonen öppnar du en dialogruta där du skapar och redigerar hyperlänkar.  
Hyperlänkdialog  
Välj vilken typ av hyperlänk du vill infoga med hjälp av symbolerna.  
Kommandoknappar  
I den här dialogrutan finns följande kommandoknappar.  
Överta  
Klicka här om du vill spara inmatningarna och stänga dialogrutan.  
Stäng  
Klicka på den här kommandoknappen om du vill lämna dialogrutan utan att spara.  
Hjälp  
Klicka på den här kommandoknappen om du vill använda hjälpen.  
Tillbaka  
Klicka här om du vill ångra inmatningarna.  
Internet  
På sidan Internet i hyperlänkdialogen kan du redigera hyperlänkar med WWW-, FTP - eller Telnet-adresser.  
Fälten Loginnamn, Lösenord och Anonym användare är bara tillgängliga för FTP-adresser.  
Typ av hyperlänk  
Internet  
Välj det här alternativet om du vill skapa en http-hyperlänk.  
FTP  
Välj det här alternativet om du vill skapa en FTP-hyperlänk.  
Telnet  
Välj det här alternativet om du vill skapa en Telnet-hyperlänk.  
Mål  
Webbläsare  
Om du klickar på den här ikonen startas webbläsaren, och med den kan du ladda en URL-adress.  
Kopiera sedan adressen till urklippet och klistra in den i fältet Mål.  
Mål i dokumentet  
Öppnar dialogrutan Mål i dokumentet.  
Där kan du välja mål i ett dokument och koppla det till mål-URL-adressen med hjälp av kommandoknappen Överta.  
Välj här till vilket ställe i måldokumentet du vill hoppa när länken aktiveras.  
Om du klickar på den här kommandoknappen, infogas målet i fältet Mål i hyperlänkdialogen.  
När hyperlänken är fullständig, klickar du på Stäng för att lämna den här dialogrutan.  
Då är länken definierad.  
Loginnamn  
För FTP-adresser kan du ange ditt loginnamn här.  
Lösenord  
För FTP-adresser kan du ange ditt lösenord här.  
Anonym användare  
Markera den här rutan om du vill logga in på FTP-adressen som anonym användare.  
Fler inställningar  
Här gör du ytterligare inställningar för den nya hyperlänken.  
Ram  
Form  
Här väljer du om hyperlänken ska skapas som text eller kommandoknapp ("Button").  
Händelser  
Genom att klicka på den här symbolen öppnar du dialogrutan Tilldela makro, där du kan förse en händelse som "Mus över objekt" eller "Utför hyperlänk "med en egen programkod.  
Text  
Skriv här den text som ska visas som läsbar text till hyperlänken eller etikett för kommandoknappen.  
Namn  
E-post & nyheter  
På sidan E-post & nyheter i dialogrutan Hyperlänk kan du redigera hyperlänkar för e-post - eller nyhetsadresser.  
E-post & nyheter  
E-post  
Med det här alternativet bestämmer du att hyperlänken hänvisar till en e-postadress.  
När du klickar på hyperlänken öppnas ett nytt meddelandedokument till mottagaren.  
Nyheter  
Med det här alternativet bestämmer du att hyperlänken hänvisar till en nyhetsadress.  
När du klickar på hyperlänken öppnas ett nytt meddelandedokument till diskussionsgruppen.  
Mottagare  
Här skriver du mottagarens fullständiga adress, i form av mailto:name@provider.com eller news:gruppe.server.com.  
Du kan också använda dra-och-släpp.  
Datakällor  
Den här kommandoknappen visar eller döljer datakällvyn.  
Angående  
Här anger du ärendet som sätts in i ärendefältet i det nya meddelandedokumentet.  
Dokument  
På sidan Dokument i hyperlänkdialogen kan du redigera hyperlänkar till valfria dokument och mål i dokumenten.  
Dokument  
Här väljer du dokument.  
Sökväg  
Öppna fil  
Den här ikonen öppnar dialogrutan Öppna fil, där du kan välja en fil.  
Mål i dokumentet  
Här väljer du målet.  
Mål  
Här kan du ange ett mål för hyperlänken i det dokument som du har angett i fältet Sökväg.  
Mål i dokumentet  
Genom att klicka här öppnar du dialogrutan Mål i dokumentet, där du kan välja ett mål bland dem som finns i dokumentet.  
URL  
Här ser du den URL-adress som är resultatet av uppgifterna i Sökväg och Mål.  
Nytt dokument  
På sidan Nytt dokument i hyperlänkdialogen kan du skapa en hyperlänk till ett nytt dokument och skapa det nya dokumentet direkt.  
Nytt dokument  
Här anger du det nya dokumentets namn, sökväg och typ.  
Redigera direkt  
Med det här alternativet skapas det nya dokumentet och laddas direkt för redigering.  
Redigera senare  
Med det här alternativet skapas det nya dokumentet som fil, men laddas inte.  
Fil  
Välj ut sökväg  
Den här symbolen öppnar dialogrutan Välj ut sökväg, där du kan välja en sökväg.  
Filtyp  
Här väljer du filtypen för det nya dokumentet som ska skapas.  
Föregående sida  
Med den ikonen hoppar du till föregående sida i dokumentet.  
Du kan bara välja den här funktionen om du har valt funktionen Förhandsgranskning på menyn Arkiv.  
Föregående sida  
Nästa sida  
Med den här ikonen hoppar du till nästa sida i dokumentet.  
Den här funktionen går bara att välja om du har valt funktionen Förhandsgranskning på Arkiv -menyn.  
Nästa sida  
Till början av dokumentet FÃ¶rsta sidan  
Genom att klicka på den här ikonen hoppar du till första sidan i dokumentet.  
Till början av dokumentet FÃ¶rsta sidan  
Till slutet av dokumentet Sista sidan  
Genom att klicka på den här ikonen hoppar du till sista sidan i dokumentet.  
Till slutet av dokumentet Sista sidan  
Förhandsgranskning  
Genom att klicka på den här kommandoknappen återvänder du till den normala dokumentvyn.  
Förhandsgranskning  
Explorer på / av  
Med den här ikonen sätter du på eller stänger av Explorer för datakällor.  
Ikonen finns på Databaslisten.  
Explorer på / av  
I Explorer för datakällor ser du datakällorna som är registrerade i %PRODUCTNAME med deras länkar, sökningar och tabeller.  
Skapa förbindelse - när du markerar en tabell eller en sökning skapas en förbindelse till datakällan.  
Tabeller och namnet på den valda sökningen eller tabellen i fetstil.  
Du måste skapa en förbindelse till datakällan innan du t.ex. kan infoga en kopierad tabell där.  
På snabbmenyn i Explorer för datakällor finns följande kommandon som är relaterade till den aktuella posten som visas inverterat:  
Kommandona på snabbmenyn skiljer sig åt beroende på om det redan finns en koppling till databasen eller inte.  
Kommandot Stäng förbindelse visas t.ex. först när det finns en koppling.  
Snabbmeny till en datakällhuvudpost  
Administrera datakällor  
Öppnar dialogrutan Administrera datakällor.  
SQL  
Öppnar dialogrutan Utför SQL-sats.  
Stäng förbindelse  
Stänger förbindelsen till datakällan.  
Se Verktyg - Alternativ - Datakällor - Förbindelser.  
Byt namn (för tabell, vy, sökning)  
När du har valt det här kommandot kan du byta namn på posten.  
Mata bara in det nya namnet.  
Du kan också dubbelklicka på posten eller markera den och trycka på F2.  
Databasen måste stödja namnbytet annars får det här kommandot ingen effekt.  
Fler kommandon på snabbmenyn till "Länkar"  
Fler kommandon på snabbmenyn till en enskild länk  
Fler kommandon på snabbmenyn till "Sökningar"  
Nytt sökningsutkast  
Öppnar fönstret Sökningsutkast.  
Mata in nytt SQL-kommando  
Med det här kommandot öppnar du sökningen om du direkt vill ange ett SQL-kommando.  
Fler kommandon på snabbmenyn till en enskild sökning  
Redigera sökning  
Med det här kommandot öppnar du sökningen i utkastvy n.  
Radera sökning  
Sökningar raderas fysiskt.  
Kopiera sökning  
Kopierar sökningen till urklippet.  
Därifrån kan du t.ex. klistra in den i ett textdokument.  
När du har valt kommandot Klistra in visas dialogrutan Infoga databaskolumner.  
Fler kommandon på snabbmenyn till "Tabeller"  
Nytt vyutkast  
Öppnar fönstret Sökningsutkast.  
Vyn utformas och används som en sökning.  
Klistra in tabell  
Klistrar in en tabell från urklippet i den markerade tabellcontainern.  
AutoPilot Kopiera tabell visas.  
Relationsutkast  
Öppnar fönstret Relationsutkast.  
Fler kommandon på snabbmenyn till en enskild tabell  
Kopiera tabell  
Kopierar den markerade tabellen till urklippet.  
Fler kommandon på snabbmenyn till en vy  
Radera vy  
Raderar den markerade vyn.  
Kopiera vy  
Kopierar den markerade vyn till urklippet.  
Klistra in vy  
Klistrar in en vy från urklippet i den markerade tabellcontainern.  
AutoPilot Kopiera tabell visas.  
Sortera stigande  
Genom att klicka på den här ikonen sorterar du data i det markerade fältet i stigande ordning.  
Data i det markerade fältet sorteras i stigande ordning när du klickar på den här ikonen.  
Textfält sorteras alfabetiskt (A-Z), numeriska fält sorteras stigande (0-9).  
Sortera stigande  
Data i det markerade fältet sorteras alltid.  
Ett datafält är markerat, när markören står i det.  
I tabeller kan du även klicka på tillhörande kolumnhuvud.  
Då öppnas en dialogruta där du kan kombinera flera sorteringskriterier.  
Sortera fallande  
Genom att klicka på den här ikonen sorterar du data i det markerade fältet i fallande ordning.  
Data i det markerade fältet sorteras i fallande ordning när du klickar på den här ikonen.  
Textfält sorteras alfabetiskt (Z-A), numeriska fält sorteras fallande (9-0).  
Sortera fallande  
AutoFilter  
AutoFilter-funktionen filtrerar dataposterna enligt innehållet i det datafält som är markerat.  
AutoFilter  
Ställ markören i det datafält, enligt vars innehåll Du vill filtrera och klicka på ikonen AutoFilter.  
Nu visas endast dataposter med samma innehåll som det markerade datafältet.  
Om Du vill att endast kunder från Göteborg ska visas i en kunddatabas så klickar Du på ett datafält med innehållet "Göteborg".  
AutoFilter filtrerar då ut samtliga kunder från Göteborg från databasen åt dig.  
Du kan upphäva det inställda AutoFiltret igen med ikonen Ta bort filter / sortering.  
Om Du vill filtrera enligt flera datafält samtidigt klickar Du på ikonen Standardfilter..., varvid en dialogruta öppnas, där Du kan kombinera flera filtreringskriterier.  
Ta bort filter / sortering  
Här upphäver du alla inställda AutoFilter eller sorteringar.  
Ta bort filter / sortering  
I sökningsutkastet ångrar du alla sökkriterier.  
Ett formulärbaserat filter raderas helt.  
Uppdatera  
Data läses in på nytt.  
Detta kan t.ex. vara lämpligt om du vill visa det aktuella databasinnehållet vid delad åtkomst till databaser i ett nätverk.  
Uppdatera  
Om du klickar länge på ikonen öppnas en undermeny med följande kommandon:  
Uppdatera - visar innehållet i databastabellen på nytt.  
Använd det här kommandot när tabellens struktur har ändrats.  
Infoga databaskolumner  
Här infogas alla fält i en markerad datapost på markörens position i det aktuella dokumentet.  
Ikonen är bara synlig om det aktuella dokumentet är ett text - eller tabelldokument.  
Det finns mer information om detta i %PRODUCTNAME Writer - resp. $[officename Calc-hjÃ¤lpen.  
Data i text  
I datakällvyn markerar du dataposten som du vill infoga i dokumentet och klickar sedan på ikonen Data i text.  
Dataposten infogas vid markörens position i dokumentet och innehållet i datapostens enskilda fält kopieras till en tabellkolumn.  
Du kan även markera flera dataposter och överföra dem till dokumentet genom att klicka på ikonen.  
Varje enskild datapost läggs då in på en ny rad.  
I datakällvyn markerar du de dataposter som du vill infoga i dokumentet och klickar sedan på ikonen Data i text.  
Då öppnas dialogrutan Infoga databaskolumner.  
Den här dialogrutan öppnas även när du drar och släpper data från en databas i datakällvyn till dokumentet eftersom du först måste ange om data ska infogas som Tabell, Fält eller Text.  
De inställningar för infogning av data som Du anger i den här dialogrutan sparas och gäller nästa gång dialogrutan öppnas.  
Denna möjlighet att spara beror på databasen och rymmer inställningar för maximalt fem databastabeller.  
Om data infogas som tabell i dokumentet sparas dock inte tabellens egenskaper.  
Samma formatmall används då automatiskt nästa gång som data infogas i tabellen om Du inte ändrar inställningarna.  
Tabell  
Här infogas de data, som är markerade i datakällvyn, som tabell i dokumentet.  
De data som har markerats infogas som tabell i dokumentet om du väljer alternativet Tabell i dialogrutan Infoga databaskolumner.  
I dialogrutan bestämmer du dessutom vilka databasfält respektive -kolumner som ska övertas och hur texttabellen ska formateras.  
Tabell  
I området Tabell väljer du med pilknapparna vilka av databastabellens kolumner som ska användas till texttabellen.  
Databaskolumner  
I den här listrutan finns alla de kolumner i databastabellen som du ännu inte har överfört till listrutan Tabell.  
Posterna står i alfabetisk ordning.  
Markera den databaskolumn vars innehåll du vill infoga i texttabellen.  
Tabell  
I listrutan Tabell visas alla databaskolumner som du har valt att infoga i dokumentet.  
Varje post tilldelas en kolumn i den tabell som ska infogas i dokumentet.  
Hur data sedan placeras i texttabellen bestäms av posternas ordningsföljd i listrutan Tabell.  
=>>  
Om du klickar på den här kommandoknappen övertas alla databasfält för att infogas i dokumentet.  
->  
Klicka på denna kommandoknapp om databasfältet som markerats i listrutan Databaskolumner ska övertas i texttabellen.  
Du kan också välja en post genom att dubbelklicka på den.  
< -  
Klicka på denna kommandoknapp om databasfältet som markerats i listrutan Tabell inte ska övertas i texttabellen.  
<<=  
Alla databasfält som skulle ha infogats i dokumentet tas bort ur listrutan Tabell om du klickar på den här kommandoknappen.  
Infoga tabellöverskrift  
Här kan du göra inställningar som gäller texttabellens överskrift.  
Infoga tabellöverskrift  
Markera den här kryssrutan om en överskriftsrad för kolumnerna ska infogas i texttabellen.  
Använd kolumnnamn  
Med detta alternativ används databastabellens fältnamn som överskrift för de enskilda kolumnerna i texttabellen.  
Skapa bara rad  
Med detta alternativ infogas en tom överskriftsrad i texttabellen.  
Du kan sedan i dokumentet definiera överskrifter som inte motsvarar databasfältens namn.  
Format  
Här kan du välja det format i vilket databasfältens innehåll ska infogas i dokumentet.  
Från databas  
Med detta alternativ övertas databasformaten.  
Urval  
I urvalslistan väljer du ett format i vilket fältinnehållet ska infogas i dokumentet.  
Nummerformaten som finns här är bara tillgängliga för vissa databasfält, t.ex. numeriska eller booleska fält.  
Om ett databasfält i textformat är markerat, kan du inte välja några format i urvalslistan eftersom textformatet bibehålls automatiskt då.  
Om det format som du vill ha inte finns med, så väljer du posten "Fler format..." för att bestämma det önskade formatet i dialogrutan Talformat.  
När ett talformat tilldelas med hjälp av urvalslistan, gäller detta alltid det databasfält som markerats i listrutan Databaskolumner.  
Om dessa data ska infogas som tabell i dokumentet och du har aktiverat det motsvarande alternativet Tabell, så kan du även välja ett databasfält i listrutan Tabell för att bestämma dess formatering.  
I det här fallet påverkar ändringen av talformatet alltid den sist markerade posten, oavsett om databasfältet har valts i listrutan Databaskolumner eller i listrutan Tabell.  
Egenskaper...  
Via den här kommandoknappen öppnar du dialogrutan Tabellformat där du kan definiera tabellens egenskaper.  
Till dessa räknas exempelvis inramningen, bakgrunden, olika justeringsalternativ och kolumnbredderna.  
AutoFormat...  
Med den här kommandoknappen öppnar du dialogrutan AutoFormat där tabellen kan formateras automatiskt.  
I den här dialogrutan kan du välja en formatmall som används direkt när tabellen infogas.  
Fält  
Välj det här alternativet om det ska infogas fältkommandon i dokumentet för de data som har markerats i datakällvyn.  
För de data som har markerats i datakällvyn infogas fältkommandon i dokumentet om du väljer alternativet Fält i dialogrutan Infoga databaskolumner.  
Dessa databasfält står sedan som platshållare för de enskilda databaskolumnerna och kan användas för standardbrev (kopplad utskrift).  
Med ikonen Data i fält anpassas fältens innehåll till den aktuella markerade dataposten.  
Ifall flera dataposter är markerade när funktionen Data i text väljs, så infogas fälten för kopplad utskrift ett motsvarande antal gånger.  
Mellan de enskilda fältkommando-blocken som ska infogas i dokumentet infogas i detta fall automatiskt ett fältkommando av typen "Nästa datapost".  
I dialogrutan Infoga databaskolumner bestämmer Du vilka databasfält som ska infogas i dokumentet och hur styckena ska formateras.  
Fält  
I området Fält väljer Du med pilknappen de av databastabellens kolumner för vilka motsvarande fältkommandon ska infogas i det aktuella dokumentet.  
Databaskolumner  
I denna listruta finns alla de kolumner i databastabellen som Du kan överta i urvalslistrutan för infogning i dokumentet.  
Posterna står i alfabetisk ordning.  
Markera den databaskolumn som Du vill använda för infogning i dokumentet.  
=>  
Klicka på denna kommandoknapp om posten som markerats i listrutan Databaskolumner ska övertas i urvalsfältet.  
Du kan också välja en post genom att dubbelklicka på den.  
Urval  
I urvalsfältet visas alla databaskolumner som Du har valt för infogning i dokumentet.  
Här kan Du även skriva in en extra text som också ska infogas.  
Hur data sedan placeras i dokumentet bestäms av posternas ordning i urvalsfältet.  
Om Du infogar en radbrytning med returtangenten, så infogas i dokumentet på detta ställe också en (stycke -) brytning.  
Styckeformatmall  
De infogade styckena formateras som standard med den aktuella styckeformatmallen.  
I listrutan Styckeformatmall motsvarar denna formatering posten "ingen".  
Här kan du vid behov välja en annan styckeformatmall som ska användas för stycket som infogas.  
I listrutan finns alla styckeformatmallar som är definierade i %PRODUCTNAME och som administreras i mallkatalogen.  
Text  
Välj det här alternativet om de data som har markerats i datakällvyn ska infogas som text i dokumentet.  
Innehållet i de data som har markerats i datakällvyn kommer att infogas som text i dokumentet om du väljer alternativet Text i dialogrutan Infoga databaskolumner.  
I dialogrutan bestämmer du vilket fältinnehåll som ska infogas i dokumentet från databasen och hur styckena ska formateras.  
Ifall flera dataposter är markerade när funktionen Data i text väljs, så infogas databasinnehållen ett motsvarande antal gånger.  
Text  
I området Text väljer Du med pilknappen för vilka av databastabellens kolumner fältinnehållen ska infogas i det aktuella dokumentet.  
Data i fält  
Här uppdateras innehållet i databasfälten med de markerade dataposterna.  
Ikonen är bara synlig om det aktuella dokumentet är ett textdokument.  
Data i fält  
Standardfilter  
Med den här ikonen filtrerar Du data enligt särskilda kriterier.  
Med funktionen AutoFilter kan Du bara filtrera efter ett enda kriterium men i den här dialogrutan kan Du kombinera flera kriterier.  
Standardfilter...  
Om Du har använt funktionen AutoFilter för att utföra en automatisk filtrering på ett markerat fält innan Du öppnar dialogrutan Filter, visas det aktiverade filtret när Du öppnar dialogrutan Filter.  
Om du samtidigt har markerat ett särskilt fält inom den filtrerade dataposten visas detta tilläggsval korrekt som en OCH-länk när dialogrutan Filter öppnas. %PRODUCTNAME tolkar ditt urval enligt mönstret "filtrerade dataposter" OCH "markering "eftersom du har valt ut en datapost bland de filtrerade dataposterna.  
Om du öppnar dialogrutan Filter visas alltså alla filter som redan används. %PRODUCTNAME känner igen en markering som du har gjort och visar den korrekta tolkningen i Filter -dialogrutan.  
När du ska utföra en ny filtrering kan du naturligtvis ändra de filtreringsvillkor som ställts in automatiskt av %PRODUCTNAME i Filter -dialogrutan.  
Du kan upphäva det inställda filtret igen med ikonen Ta bort filter / sortering.  
Standardfilter / filter  
I den här dialogrutan anger Du logiska villkor för filtrering av data i en tabell.  
I tabelldokument heter dialogrutan Standardfilter och i databastabeller eller -formulär heter den Filter.  
Dialogrutan Filter innehåller inte kommandoknappen Fler.  
Filterkriterier  
Ett standardfilter kan Du definiera genom att ange länktyp, fältnamn, logiskt villkor och ett värde respektive en kombination av argument.  
Operator  
För efterföljande argument kan Du välja mellan de logiska operatorerna OCH och ELLER.  
Fältnamn  
Välj i listrutan det fältnamn som Du vill föra in i argumentet i den aktuella tabellen.  
Om det inte finns någon text som anger fältnamnet visas i stället kolumnbeteckningen här.  
Villkor  
I listrutan kan Du välja mellan flera jämförelseoperatorer med vilka posterna i fälten Fältnamn och Värde ska länkas.  
Värde  
Här anger Du det värde enligt vilket fältet ska filtreras.  
I %PRODUCTNAME Calc-tabeller visas i ett listfält alla möjliga värden som kan föras in i kolumnen Fältnamn.  
Här kan Du också välja posterna "tom" och "inte tom "för att kunna filtrera mellan tomma respektive ifyllda poster.  
Om Du använder filterfunktionen i databastabeller eller -formulär, anger Du i textfältet ett värde som ska användas för filtrering.  
Fler>>  
Jämförelseoperatorer  
I dialogrutan Standardfilter kan Du under Villkor välja följande jämförelseoperatorer:  
Jämförelseoperator  
Effekt  
Lika med (=)  
Visar de värden som är lika med villkoret.  
Mindre än (<)  
Visar de värden som är mindre än villkoret.  
Större än (>)  
Visar de värden som är större än villkoret.  
Mindre än eller lika med (< =)  
Visar de värden som är mindre än eller lika med villkoret.  
Större än eller lika med (> =)  
Visar de värden som är större än eller lika med villkoret.  
Inte lika med (< >)  
Visar de värden som inte är lika med villkoret.  
största  
Visar de N (numeriskt värde som parameter) största värdena.  
minsta  
Visar de N (numeriskt värde som parameter) minsta värdena.  
största%  
Visar de största N% (numeriskt värde som parameter) av det totala antalet värden.  
minsta%  
Visar de minsta N% (numeriskt värde som parameter) av det totala antalet värden.  
Sortera  
Sortera  
Sortering  
Här kan Du ange sorteringskriterier för hur data ska visas.  
Med funktionerna Sortera stigande och Sortera fallande kan Du bara sortera enligt ett enda kriterium, men i den här dialogrutan kan Du kombinera flera kriterier.  
Du kan upphäva en utförd sortering genom att klicka på ikonen Ta bort filter / sortering.  
Sortering  
Här anger Du sorteringskriterierna.  
Om Du därefter anger ytterligare sorteringskriterier så sorteras de data som överensstämmer med det överordnade kriteriet enligt nästa kriterium.  
För varje förnamn sorteras sedan dataposterna fallande efter efternamn.  
Fältnamn  
Här väljer Du namnet på det datafält, efter vars innehåll sorteringen ska ske.  
Ordning  
Här anger Du om sorteringen ska ske i stigande eller fallande ordning.  
därefter  
Ange ytterligare underordnade sorteringskriterier i de övriga fälten.  
Sök datapost  
Med den här ikonen kan du söka efter bestämda värden i datafält.  
I formulär och databastabeller kan du söka efter särskilda värden i datafält, listrutor och kryssrutor.  
Vid sökning i en tabell genomsöks datafälten i den aktuella tabellen.  
Vid sökning i ett formulär genomsöks de datafält i tabellen som är länkade till formuläret.  
Den sökning som beskrivs här utförs av din programversion av %PRODUCTNAME Base.  
Om du vill använda SQL-servern för en sökning i en databas använder du ikonen Formulärbaserat filter på Formulärlisten.  
Det går även att använda sökfunktionen för tabellkontrollfält.  
Om du använder sökfunktionen för ett markerat tabellkontrollfält, kan du söka i de enskilda kolumnerna i tabellkontrollfältet som motsvarar databaskolumnerna i den länkade databastabellen.  
Sök efter  
Här väljer du vad du vill söka efter.  
Text:  
Skriv sökordet i kombinationsfältet eller välj det i listan.  
Om markören står i ett fält när dialogrutan öppnas och fältet innehåller enbart text (utan tabbar och radbrytningar), införs den här posten automatiskt i kombinationsfältet i sökdialogrutan.  
Ändra posten men tänk på att tabbar och radbrytningar inte kan bearbetas vid sökning i ett formulär.  
Alla sökord under en session sparas så länge tabellen eller formulärdokumentet är öppet.  
Om du har gjort flera sökningar och skulle vilja använda ett tidigare använt sökord igen, kan du hitta det i listrutan.  
Fältinnehållet är NULL  
Om det här alternativet är markerat, görs sökningen efter fält som saknar innehåll.  
Fältinnehållet är inte NULL  
Med det här alternativet hittas fält som har innehåll.  
Område  
Här bestämmer du i vilka fält sökningen ska göras.  
Formulär  
Här kan du ange i vilket logiskt formulär sökningen ska göras.  
Det här kombinationsfältet visas bara om det aktuella dokumentet är ett formulärdokument med mer än ett logiskt formulär.  
Det visas alltså inte vid sökning i tabeller eller sökningar.  
Ett formulärdokument kan innehålla flera logiska formulär.  
De utgörs av enskilda formulärkomponenter som alltid är länkade till en tabell.  
Antag att Du har ett formulär (som hänför sig till Tabell A) med ett underformulär (som hänför sig till Tabell B).  
Ett överordnat och ett underordnat formulär är alltid logiska formulär.  
Ditt formulärdokument består alltså av två logiska formulär.  
Kombinationsfältet innehåller namnen på alla logiska formulär för vilka det finns kontrollfält.  
Det logiska formulär vars kontrollfält var markerat när du öppnade dialogrutan är förinställt.  
Alla fält  
Aktivera det här alternativet om sökningen ska göras i alla fält.  
Vid sökning i formulär genomsöks alla fält i det logiska formulär som har ställts in under Formulär.  
Vid sökning i tabellkontrollfältet genomsöks alla kolumner som är länkade till ett giltigt datafält i en databastabell.  
Fälten i det aktuella logiska formuläret behöver inte vara identiska med fälten i formulärdokumentet.  
Om formulärdokumentet innehåller fält som hänvisar till flera datakällor (alltså flera logiska formulär), leder alternativet Alla fält till att bara de fält i formulärdokumentet genomsöks som är länkade till en datakälla.  
Enskilt fält  
Om du väljer det här alternativet, kan du ange ett datafält som ska genomsökas.  
Inställningar  
Här kan du göra olika inställningar av sökningen.  
Position  
Ange här på vilket sätt sökordet förhåller sig till fältinnehållet.  
Följande möjligheter finns:  
var Du vill i fältet  
Alla fält hittas som innehåller sökbegreppet någonstans: i början, i slutet eller däremellan.  
i fältets början  
Alla fält hittas som inleds med sökbegreppet.  
Vid fältslut  
Alla fält hittas som avslutas med sökbegreppet.  
i hela fältet  
Alla fält hittas där innehållet enbart utgörs av (hela) sökbegreppet.  
Om rutan Platshållaruttryck är markerad är den här funktionen inte tillgänglig.  
Använd fältformatering  
Om den här rutan är markerad, tas vid sökningen hänsyn till fältformateringarna i det aktuella dokumentet.  
Fältformateringar är alla synliga formateringar som kan ställas in med följande alternativ:  
i tabellutkast vid fältegenskaperna,  
i datavyn över kolumnformateringen,  
i formuläret över kontrollfältegenskaperna.  
Om du vill söka i data i datavyn över en tabell eller i ett formulär, kan du välja om sökningen ska ta hänsyn till den för tillfället synliga formateringen eller till en standardformatering i databasen.  
Om rutan inte är markerad görs sökningen i databasen med den formatering som är sparad där.  
Exempel:  
Anta att Du har ett datumfält som har sparats med formatet "DD.MM.ÅÅ" (t ex 17.02.65) i databasen.  
Välj t ex formatet "DD MMM ÅÅÅÅ" för datavyn, så att datumet visas så här: "17 feb 1965 ".  
Efter en sådan fältformatering hittas en datapost som innehåller datumet 17 februari bara med följande inställningar:  
Använd fältformatering  
Sökord  
på  
"feb" hittas, däremot inte "2 ".  
av  
"2" hittas, däremot inte "feb ".  
Du bör göra sökningen med fältformatering, eftersom den i annat fall utgår från (interna) standardformateringar, vilket kan leda till oönskade resultat.  
Följande exempel visar vilka problem som kan uppstå om Du söker utan fältformatering.  
De beror av vilken databas som används och inträffar bara vid vissa interna standardformateringar:  
Sökresultat  
Orsak  
"5" hittar klockslaget "14:00:00 "  
Tidfält är inte definierade i dBase-databaser och måste simuleras.  
För intern representation av klockslaget "14:00:00" används 5.  
Med "00:00:00" hittas alla dataposter i ett rent datumfält  
Internt sparar databasen ett datumvärde i ett kombinerat datum - och tidfält.  
"45,79" hittar inte "45,79 "trots att alternativet hela fältet har valts under Position.  
Den synliga representationen motsvarar inte den interna lagringen.  
Om värdet 45,789 t ex har införts i ett fält av typen Tal / Dubbelt i databasen, och formateringen för visning är inställd så att bara två decimaler visas, hittas "45,79" bara i en sökningen med fältformatering.  
Standardformateringarna är i det här fallet sådana som hänför sig till den interna lagringen av data.  
För Dig som användare är de inte alltid så lätta att känna igen - särskilt inte när de används för att simulera datatyper (t ex när det gäller tidsfält i dBase-databaser).  
I det enskilda fallet beror detta på vilken databas och datatyp som används.  
Tänk på att Du vid en sökning med fältformatering alltid är på den säkra sidan om Du bara vill hitta data av den typ som Du ser på skärmen.  
Detta gäller särskilt fält av typen datum, klockslag, datum / klockslag eller tal / dubbel.  
En sökning utan fältformatering kan dock vara att föredra, eftersom den går mycket snabbare.  
Därför kan det vara bra att välja detta alternativ för stora datauppsättningar där inga formateringsproblem föreligger.  
Om du söker "med fältformatering" i kryssrutor, får du resultatet "1 "för markerade rutor, för omarkerade "0" och för obestämda (gråtonade) en tom sträng.  
Om sökningen görs utan Använd fältformatering, får du de språkberoende standardvärdena "SANN" eller "FALSK ".  
Vid sökning i listfält "med fältformatering" hittas de texter som visas i listrutorna, och vid sökning "utan fältformatering "hittas de innehåll som motsvarar den normala fältformateringen.  
Exakt sökning  
Vid exakt sökning tas hänsyn till versaler och gemener.  
Sök bakåt  
Här kan du vända sökriktningen.  
I annat fall görs sökningen framåt (från den första dataposten till den sista).  
Från början / slutet  
Om den här rutan är markerad, startas sökningen på nytt.  
Vid en framåtsökning (när kryssrutan Sök bakåt inte är markerad) börjar sökningen om med den första dataposten i tabellen; vid en bakåtsökning (när kryssrutan Sök bakåt är markerad) med den sista dataposten.  
Markera den här rutan om du inte vill gå vidare med en sökning utan upprepa den.  
När en sökning påbörjas startar den alltid med den första eller sista dataposten.  
Jokerteckenuttryck  
Markera den här rutan om du vill söka med ett jokertecken (* eller?).  
Markera den här rutan om sökordet innehåller ett jokertecken.  
Följande jokertecken tillåts:  
Jokertecken  
Betydelse  
Exempel  
?  
för exakt ett valfritt tecken  
"?ök" hittar "sök", "kök", "rök "osv  
"J?nsson" hittar t.ex. "Jansson", "Jonsson "och "Jönsson".  
*  
för 0 eller flera valfria tecken  
"*-*" hittar "ZIP-drive "och "cd-rom"  
"J*son" hittar alla poster som börjar med "J "och slutar med "son" (t.ex. Jansson, Johansson, Josefson).  
Om jokertecknet "?" eller "* "själv ska utgöra ett tecken i sökordet, ska det föregås av ett omvänt snedstreck, alltså "\?" respektive "\* "(utan citattecknen).  
Men det behövs bara när du gör en sökning med jokertecken.  
I "normalt" läge behandlas jokertecknen som vanliga tecken.  
Reguljärt uttryck  
Om du markerar den här rutan kan du söka med reguljära uttryck.  
I reguljära uttryck används särskilda tecken som styr sökförloppet.  
Det kan röra sig om jokertecken och tecken som definierar en viss sökning.  
Du kan använda samma reguljära uttryck som i dialogrutan Sök och ersätt i %PRODUCTNAME.  
Den senare typen är dock ofta tillräcklig vid normal användning och enklare att hantera.  
Om du använder sökning efter reguljära uttryck motsvaras sökning med jokertecken av följande tecken:  
Sökning med jokertecken  
Sökning efter reguljära uttryck  
?  
.  
*  
.*  
Status  
På statusraden visas den aktuella dataposten i sökresultatet.  
Om sökningen har nått slutet (respektive början) på tabellen, fortsätter den automatiskt från början (respektive slutet).  
Alltefter sökriktning visas då motsvarande upplysning.  
För mycket stora datauppsättningar kan förmedlingen av dataposter ta lite tid vid sökning i omvänd sökriktning.  
Du får då information på statusraden om att dataposterna fortfarande håller på att genomsökas.  
Sök / Avbryt  
Med den här kommandoknappen startar respektive avbryter Du sökningen.  
Med kommandoknappen Sök startar Du sökningen.  
Om den gav resultat, markeras det funna datafältet med en röd rektangel.  
Du kan därefter fortsätta sökningen med Sök eller upprepa den med inställningen Från början respektive Från slutet.  
En pågående sökning kan Du avbryta genom att åter klicka på samma kommandoknapp.  
Om Du vill avsluta sökningen och stänga dialogrutan klickar Du på Stäng.  
Stäng  
Inställningarna för den senaste sökningen sparas tills Du avslutar %PRODUCTNAME.  
Om Du har flera tabeller eller formulär öppna, kan Du ställa in ett separat sökalternativ för vart och ett av dem.  
Om Du sedan stänger dokumenten ett och ett, sparas sökalternativen i det sista.  
Formulärbaserat filter  
Med den här ikonen ser Du till att databasservern filtrerar data i ett formulär enligt bestämda kriterier.  
Med ett formulärbaserat filter kan Du söka snabbare (eftersom det som regel är en snabbare databasserver som utför sökningen) och definiera mer komplexa sökvillkor än vad som är fallet i normala sökningar, som Du startar på formulärlisten med t ex ikonen Sök datapost....  
Formulärbaserat filter  
Använd filter  
Här växlar du mellan filtrerad och ofiltrerad vy av formuläret.  
Om ikonen är intryckt visas den filtrerade vyn, annars visas den ofiltrerade.  
Om ikonen är gråtonad har inget filter definierats.  
Använd filter  
Med den här funktionen sparar du ett formulärbaserat filter så att du sedan inte behöver definiera det på nytt.  
Datakälla som tabell  
Här aktiverar och inaktiverar du tabellvyn i formulärvyn.  
Om ikonen är intryckt visas tabellen i en ram i övre kanten av formuläret, annars visas bara formuläret.  
Datakälla som tabell  
I den gemensamma vyn är tabellen och formuläret i många avseenden likställda.  
Det betyder att en datapost som Du markerar i tabellen genast visas i formuläret, och att en ändring i formuläret också visas i tabellen (och omvänt).  
Tabellen kan aldrig visa mer än ett logiskt formulär även om dokumentet innehåller flera.  
Du kan flytta ramkanten på tabellvyn med musen.  
Om Du håller ner Ctrl-tangenten och dubbelklickar på ett tomt område i den förankrade ramen, förvandlas den till ett fritt fönster.  
Om Du dubbelklickar på samma sätt en gång till förankras ramen till sin senaste position.  
Den här uppdelningen av vyn i formulär och tabell kan Du även göra om Du med hjälp av utrullningslisten Formulärfunktioner har skapat ett eget formulär baserat på ett text-, tabell - eller presentationsdokument.  
Då visas t ex varje grupp av alternativfält i formuläret som en listruta i tabellvyn.  
Aktuell dokumentdatakälla  
Här visar du i datakällvyn den tabell som är kopplad till det aktuella elementet.  
Aktuell dokumentdatakälla  
Med Redigera - Byt databas kan du välja en annan tabell.  
Ställa in tabbar  
Ställ in tabbarna för det aktuella stycket eller för alla markerade stycken genom att klicka med musen på linjalen.  
I den horisontella linjalen är standardtabbarna förinställda på 2 cm avstånd mellan varandra.  
Så snart du definierar en egen tabulator står bara standardtabbarna till höger om den kvar.  
Definiera indrag, marginaler och kolumner  
Du kan definiera indrag och marginaler för aktuellt stycke, eller alla markerade stycken, med musen.  
Om Du delat in en sida i spalter, eller om markören står i en flerspaltig textram, kan Du ändra spaltbredden och mellanrummet mellan spalterna fritt genom att dra med musen på linjallisten.  
Då kan Du ändra det genom att dra med musen på linjallisten.  
Om markören står i en tabellcell kan Du på linjallisten både ändra indraget för cellens innehåll och dra i begränsningslinjerna för att ändra tabellkolumnernas indelning.  
De här symbolerna visar vänstra indraget för första raden i aktuellt stycke (övre triangeln) och vänstra indraget för övriga rader i stycket (nedre triangeln).  
Symbolen till höger på linjallisten visar höger indrag för det aktuella stycket.  
Om Du vill  
Gör Du så här  
Göra indrag från vänster  
Dra den vänstra undre markeringen åt höger med nedtryck musknapp  
Göra förstaradsindrag från vänster  
Dra den vänstra övre markeringen åt höger med nedtryckt musknapp  
Göra indrag från höger  
Dra markeringen vid högra kanten åt vänster med nedtryckt musknapp  
Om Du endast vill ändra det vänstra indraget fr o m andra raden i ett stycke håller Du Kommando Ctrl -tangenten nedtryckt och klickar på den vänstra nedre triangeln och drar den åt höger med musen.  
Eventuella tabbar i ett stycke ändras inte när Du gör ett indrag.  
Om några tabbar hamnar utanför styckemarginalerna syns de inte, men tas inte bort.  
Utför  
Visa sökresultatet genom att klicka på den här ikonen.  
Klicka på ikonen Utför så utförs SQL-sökningen och sökresultatet visas.  
Sökningen sparas dock inte.  
Den här funktionen är användbar om du t.ex. vill kontrollera sökningen igen och eventuellt ändra den.  
När du till slut sparar sökningen placeras den under fliken Sökning.  
Utför  
Radera sökning  
Om du klickar på den här ikonen, raderas sökningen och samtliga tabeller tas bort från utkastfönstret.  
Radera sökning  
Lägg till tabeller  
Välj de tabeller som ska läggas till i Utkast-fönstret genom att klicka här.  
I den här dialogrutan väljer Du de tabeller som Du vill arbeta med.  
När Du skapar en sökning eller ny tabellvy är det här som Du väljer vilka tabeller som ska ingå i sökningen respektive tabellvyn.  
För en relationsdatabas anger Du vilka tabeller som ska ställas i relation till varandra.  
Du lägger till tabeller i sökningsutkastet eller i relationsfönstret, där de visas som egna fönster med en lista över de datafält som ingår i tabellen.  
De här fönstren kan Du ändra storlek på och flytta om.  
Tabell  
Här väljer Du en tabell.  
Tabellnamn  
Klicka på namnet på den tabell som Du vill lägga till och sedan på Lägg till.  
Du kan även dubbelklicka på tabellnamnet.  
Då visas ett fönster med tabellens datafält överst i sökningsutkastet respektive relationsfönstret.  
Lägg till  
Lägg till den markerade tabellen i utkastet genom att klicka.  
Stäng  
Efter det att Du har angett vilka tabeller som Du ska arbeta med, stänger Du dialogrutan genom att klicka på den här kommandoknappen.  
Sätt på / stäng av designvy  
Om den här ikonen är intryckt visas designvyn av sökningen.  
Om den inte är intryckt visas SQL-vyn.  
Sätt på / stäng av designvy  
Utför SQL-kommando direkt  
I Native SQL-läge anger du SQL-kommandon som inte tolkas av %PRODUCTNAME utan skickas vidare direkt till datakällan.  
Om ändringarna inte kan visas i designvyn går det att växla tillbaka till designvyn.  
När det gäller Native SQL överförs SQL-strängen direkt till databassystemet utan att först utvärderas av %PRODUCTNAME.  
Om Du t ex använder ODBC-gränssnittet för databasåtkomst överlämnas SQL-strängen till ODBC-drivrutinen som därefter bearbetar den.  
Utför SQL-kommando direkt  
I normalläget är ändringarna i sökningsutkastet synkroniserade med de tillåtna ändringarna per SQL.  
Funktioner  
Om den här ikonen är intryckt, visas raden "Funktion" i nedre delen av sökningsutkastet.  
Funktioner  
Tabellnamn  
Om den här ikonen är intryckt, visas raden "Tabell" i nedre delen av sökningsutkastet.  
Tabellnamn  
Aliasnamn  
Om den här ikonen är intryckt, visas raden "Alias" i nedre delen av sökningsutkastet.  
Aliasnamn  
Entydiga värden  
Om den här ikonen är intryckt, utökas Select-satsen i SQL-sökningen i den aktuella kolumnen med parametern DISTINCT.  
Det innebär att om samma värde förekommer flera gånger kommer det bara att förtecknas en gång.  
Entydiga värden  
Urval  
Ikonen med pilen är urvalsverktyget.  
Klicka på den om du t.ex. vill återgå till det normala urvalsläget från ritläget.  
Urval  
Med den här ikonen växlar Du till det normala urvalsläget.  
I det här läget kan du markera objekt genom att klicka på dem.  
Om du samtidigt håller ner Kommando Ctrl och Skifttangenten kan du lätt ändra objektgrupperingar.  
Håll ner en tangent och klicka på flera objekt efter varandra för att markera dem gemensamt.  
Om du klickar på ett markerat objekt igen (och samtidigt fortsätter att hålla ner skifttangenten) upphävs markeringen för det här objektet.  
Objekten som är sammanfogade på det här sättet kan sedan definieras som Gruppering vilket innebär att de omvandlas till ett enda objekt.  
Om du vill redigera enskilda element i en gruppering kan du hålla ner Kommando Ctrl -tangenten, klicka med musen och på så sätt lösa enskilda objekt från grupperingen utan att gå in i den med motsvarande menykommando.  
Det går att redigera eller placera om bara vissa objekt i grupperingen.  
Då kan du markera enskilda objekt genom att dubbelklicka.  
Genom att kombinera de beskrivna metoderna kan du lätt ändra flera grupperingar och deras objekt, samt förbindelserna mellan grupperingarna.  
Med det här verktyget kan du skapa en rektangulär ram runt flera objekt.  
Alla objekt, vars omgivande rektangel ligger helt inom ramen, markeras.  
I det här läget kan du markera objekt genom att klicka på dem.  
Om du samtidigt håller ner Kommando Ctrl och Skifttangenten kan du lätt ändra objektgrupperingar.  
Håll ner skifttangenten och klicka på flera objekt efter varandra för att markera dem gemensamt.  
Om du klickar på ett markerat objekt igen (och samtidigt fortsätter att hålla ner skifttangenten) upphävs markeringen för det här objektet.  
Objekten som är sammanfogade på det här sättet kan sedan definieras som Gruppering vilket innebär att de omvandlas till ett enda objekt.  
Om du vill redigera enskilda element i en gruppering kan du hålla ner Kommando Ctrl -tangenten, klicka med musen och på så sätt lösa enskilda objekt från grupperingen utan att gå in i den med motsvarande menykommando.  
Det går att redigera eller placera om bara vissa objekt i grupperingen.  
Då kan du markera enskilda objekt genom att dubbelklicka.  
Genom att kombinera de beskrivna metoderna kan du lätt ändra flera grupperingar och deras objekt, samt förbindelserna mellan grupperingarna.  
Med det här verktyget kan Du skapa en rektangulär ram runt flera objekt.  
Alla objekt, vars omgivande rektangel ligger helt inom ramen, markeras.  
Du kan skapa en rektangulär ram och redigera det område som du definierar på detta sätt oberoende av den övriga bildytan.  
Infoga objekt Infoga objekt  
Den här ikonen öppnar utrullningslisten Infoga objekt med funktioner för infogning av objekt.  
Du kan nu med en kort klickning aktivera funktionen på nytt.  
Med en längre klickning öppnar du i stället utrullningslisten, så att du kan välja en annan funktion.  
Ikon på verktygslisten:  
Infoga objekt Infoga objekt  
När Du för första gången har valt en funktion på utrullningslisten, visas alltid ikonen för den senast infogade funktionen.  
Om Du drar bort den från verktygslisten, får Du tillbaka listen med dess olika funktioner.  
Infoga diagram  
%PRODUCTNAME Infoga %PRODUCTNAME Math-objekt Infoga formel  
Infoga ramteknik  
Infoga andra objekt  
Infoga plug-in  
Infoga applet  
AutoRättstavning  
AutoRättstavning  
HTML-källtext  
Med kommandot HTML-källtext växlar du till ett läge där du kan se HTML-sidors källtext.  
Det här kommandot visas bara när ett HTML-dokument är öppet.  
Innan du kan ställa om ett nytt dokument till HTML-källtext måste det sparas som webbsida (HTML).  
I HTML-källtextläge visas taggarna i HTML-språket.  
Du kan redigera dessa och spara dokumentet som rent textdokument.  
Ge dokumentet filnamnstillägget .html eller .htm för att markera att det är ett HTML-dokument.  
Kommandot HTML-källtext finns även på HTML-dokumentets snabbmeny när HTML-källtexten visas.  
Genom att klicka på kommandot återgår du till normalvyn igen.  
Aktuell sidformatmall  
I det här fältet på statuslisten ser du vilken sidformatmall som används.  
Om du vill redigera den, dubbelklickar du här; och om du vill byta ut den högerklickar du.  
Om du dubbelklickar på det här fältet öppnas en dialogruta där du kan redigera sidformatmallen.  
På snabbmenyn till det här fältet kan du tilldela den aktuella sidan någon av de sidformatmallar som finns i Stylist.  
Om du dubbelklickar på det här fältet öppnas en dialogruta där du kan redigera sidformatmallen.  
Om du dubbelklickar i det här fältet öppnas dialogrutan Sidformatmall, där du kan välja mall för den aktuella sidan.  
Här kan du välja ett annat pappersformat eller en annan bakgrund.  
Om du dubbelklickar i det här fältet öppnas dialogrutan Sidformatmall, där du kan välja mall för den aktuella sidan.  
Här kan du välja ett annat pappersformat eller en annan bakgrund.  
Skala  
Här ser du och kan ändra den aktuella skalan för sidvisningen.  
Om du dubbelklickar i det här fältet öppnas dialogrutan Skala, där du kan ställa in skalan.  
Om du öppnar snabbmenyn i det här fältet, får du upp en lista över de alternativa förstoringar av vyn som du kan välja bland.  
Infogningsläge  
I det här fältet visas det aktuella infogningsläget.  
Här kan du byta mellan INFGA = infoga; ÖVER = skriva över.  
Fältet är bara aktivt när markören står på formellistens inmatningsrad eller i en cell.  
Med en enkel musklickning i fältet ändrar Du läget i tur och ordning mellan de tillgängliga alternativen (utom i %PRODUCTNAME Basic-IDE, där bara tangenten Insert kan användas).  
Du kan ändra läget även med tangenten Insert när markören står i dokumentet.  
Läge:  
Effekt:  
INFGA  
I infogningsläget infogas nya tecken vid markörens position, och efterföljande text flyttas åt höger.  
Markören visas som ett lodrätt streck.  
ÖVER  
I överskrivningsläget skriver nya tecken över de som redan finns.  
Markören visas som block.  
Markeringsläge  
Här visas det aktuella markeringsläget.  
Du kan växla mellan STD = standard, UTV = utvidga och TLF = tillfoga här.  
Varje gång som du klickar i det här fältet växlar du till nästa läge.  
Visning:  
Läge:  
Effekt:  
STD  
Normalläge  
När du klickar i texten placeras textmarkören där; om du klickar på en cell gör du den till aktuell cell.  
En befintlig markering upphävs.  
UTV  
Utvidgningsläge  
Genom att klicka i texten utökar eller minskar du den aktuella markeringen till det ställe där du klickar.  
Om du klickar före eller efter den tidigare markeringen, sträcker sig den nya markeringen till början respektive från slutet av denna.  
TLF  
Kompletteringsläge  
Om du gör en ny markering finns de tidigare markeringarna kvar.  
Det uppstår en multimarkering, d.v.s. en markering som inte kan bestå av icke sammanhängande delar.  
Dokumentändring  
Om dokumentet innehåller ändringar som ännu inte har sparats, visas detta i statuslisten med en asterisk (*) i det här fältet.  
Detta gäller även för nya dokument, som ännu inte har sparats.  
Kombinerad visning  
Här visas aktuellt datum och klockslag.  
Klockslag  
I detta fält visas det aktuella klockslaget.  
Datum  
I detta fält visas det aktuella datumet.  
Klockslag  
I detta fält visar %PRODUCTNAME aktuellt klockslag.  
Storlek  
Här visas sammanfattande information om de enheter, mappar och filer som visas.  
Filter  
Med filterverktyget på grafikobjektlisten öppnar du fönstret Filter, där du kan använda filter för det markerade grafikobjeket.  
Filter  
Invertera  
Det här filtret inverterar färgvärdena i en färgbild eller värdena för ljusstyrkan i en bild i gråskalor eller svartvitt.  
Invertera  
Utjämna  
Det här filtret utjämnar kontrasterna i bilden.  
Utjämna  
Skärpa  
Det här filtret ökar kontrasterna i bilden.  
Skärpa  
Ta bort brus  
Det här filtret tar bort enstaka pixel från bilden.  
Ta bort brus  
Solarisering  
Om du klickar på den här ikonen öppnas en dialogruta där du kan ställa in solarisationen.  
Med solarisation menas en effekt som kan uppstå när fotomaterial överexponeras under framkallningen.  
Solarisationen förvränger färgerna genom att delvis invertera dem.  
Solarisering  
Parametrar  
Här ställer du in grad och typ av solarisering.  
Tröskelvärde  
I det här rotationsfältet anger du graden av ljusstyrka i procent från vilken pixlarna ska solariseras.  
Invertera  
Markera den här rutan om pixlarna som ska solariseras samtidigt ska få inverterade färger.  
Åldrande  
Om du klickar på den här ikonen öppnas en dialogruta där du kan ställa in funktionen åldrande.  
Bilden blir lite mörkare för varje gång den här funktionen aktiveras, färgerna kan ändras i riktning grått och / eller brunt.  
Åldra  
Åldringsgrad  
I det här rotationsfältet ställer du in intensiteten för åldringsgraden i%.  
Ju högre värde du väljer desto mer åldras din bild.  
Poster  
Om du klickar på den här ikonen öppnas en dialogruta där du kan definiera antalet posterfärger.  
Den här effekten baserar på reducering av färgantalet.  
På så sätt kan du få fotolika bilder att se ut som om de vara målade.  
Poster  
Posterfärger  
I det här fältet väljer du antalet färgnivåer som bilden ska reduceras till.  
Klicka sedan på OK så reduceras bilden till det här antalet färgnivåer.  
Popkonst  
Om du klickar på den här ikonen omvandlas ditt grafikobjekt till ett popkonstdokument.  
Genom färgförändring får ditt grafikobjekt en helt annan karaktär.  
Den här funktionen kan användas både på hela grafikobjektet och för ett markerat område.  
Popkonst  
Kolteckning  
Med det här kommandot visas grafikobjektet som kolteckning.  
Grafikobjektets konturer fylls i med svart och de ursprungliga färgerna undertrycks.  
Den här funktionen kan både användas för hela grafikobjektet och för ett markerat område.  
Kolteckning  
Relief  
Om du klickar på den här ikonen öppnas en dialogruta för reliefutformning.  
Här väljer du den tänkta platsen för en imaginär ljuskälla.  
Den här ljuskällan bestämmer hur skuggan faller och därmed utseendet på ett grafikobjekt som omvandlas till en relief.  
Den här funktionen kan både användas på hela grafikobjektet och för ett markerat område.  
Relief  
Ljuskälla  
I det här fältet klickar du på platsen där du vill att ljuskällan ska placeras.  
Den symboliseras av en punkt.  
Mosaik  
Med den här funktionen sammanfogas små pixelgrupper till rektangulära ytor med samma färg.  
Ju större de enskilda rektanglarna är desto detaljfattigare blir grafikobjektet.  
Mosaik  
Elementupplösning  
Bestäm här hur många pixlar som ska sammanfogas till rektanglar.  
Bredd  
Definiera bredden på de enskilda kakelplattorna med det här rotationsfältet.  
Höjd  
Definiera höjden på de enskilda kakelplattorna med det här rotationsfältet.  
Framhäv kanter  
Om du markerar den här rutan framhävs kanterna på objektet (görs skarpare).  
Grafikläge  
I listrutan Grafikläge väljer du ett visningsattribut för det markerade grafikobjektet.  
Grafikobjekt som är inbäddat eller länkat i den aktuella filen förändras inte, bara visningen av objektet ändras.  
Grafikläge  
Standard  
Visningen av grafikobjektet förändras inte.  
Gråskalor  
Ett grafikobjekt i färg visas monokromt, först i gråskalor.  
Du kan dessutom få en färgad toning av gråskalorna genom att öka värdet på en av färgregulatorerna.  
Svartvitt  
Ett grafikobjekt visas i svartvitt.  
Alla ljusstyrkevärden under 50% blir svarta, alla över 50% blir vita.  
Vattenmärke  
Grafikobjektet visas med förminskad ljusstyrka och kontrast, vilket gör att det lämpar sig som vattenmärke i bakgrunden.  
Andel rött  
I rotationsfältet Andel rött ökar eller minskar du andelen röd RGB-färgkomponent i visningen av det markerade grafikobjektet.  
Du kan välja värden från -100% (inget rött alls) till +100% (fullt värde).  
Andel rött  
Andel grönt  
I rotationsfältet Andel grönt ökar eller minskar du andelen grön RGB-färgkomponent i visningen av det markerade grafikobjektet.  
Du kan välja värden från -100% (inget grönt alls) till +100% (fullt värde).  
Andel grönt  
Andel blått  
I rotationsfältet Andel blått ökar eller minskar du andelen blå RGB-färgkomponent i visningen av det markerade grafikobjektet.  
Du kan välja värden från -100% (inget blått alls) till +100% (fullt värde).  
Andel blått  
Ljusstyrka  
I det här rotationsfältet väljer du högre eller lägre ljusstyrka i visningen av det markerade grafikobjektet.  
Du kan välja värden från -100% (bara svart) till +100% (bara vitt).  
Ljusstyrka  
Kontrast  
I rotationsfältet Kontrast ställer du in högre eller lägre kontrast i vyn över markerade grafikobjekt.  
Möjliga värden är från -100% (ingen kontrast alls) till +100% (full kontrast).  
Kontrast  
Gamma  
Här ökar eller minskar du gammavärdet för visningen av det markerade grafikobjektet.  
Du kan välja värden från 0,10 (minimal gamma) till 10 (maximal gamma).  
När ett gammavärde ändras sker en icke-linjär förändring av ljusstyrkan.  
Gamma  
Transparens  
I rotationsfältet Transparens ökar eller minskar du transparensen för visningen av det markerade grafikobjektet.  
Du kan välja värden från 0% (inte genomskinlig) till +100% (helt genomskinlig).  
Transparens  
Beskära  
Om du klickar på den här ikonen öppnas en dialogruta där du kan beskära pixelgrafik.  
Funktionen är bara tillgänglig för ett markerat pixelgrafikobjekt.  
beskära  
Allmänna kortkommandon i %PRODUCTNAME  
Här är standard-tangentkombinationerna listade som används i hela %PRODUCTNAME.  
Utföra kommando direkt med hjälp av tangentkombinationer  
Du kan starta ett stort antal funktioner i ditt program via tangentkombinationer.  
Bredvid Öppna på menyn Arkiv står exempelvis tangentkombinationen Kommando+O Ctrl+O.  
Om du vill starta funktionen via tangentkombinationen håller du ner Kommando Ctrl -tangenten och trycker på tangenten O.  
Släpp därefter båda tangenterna.  
Du kan välja mellan att använda musen eller tangentbordet för nästan alla funktioner.  
Öppna menyer direkt med hjälp av tangentkombinationer  
På menylisten är många tecken understrukna.  
Du öppnar de här menyerna genom att trycka på det understrukna tecknet och samtidigt hålla ner Alt-tangenten.  
På menyn som öppnas hittar du fler understrukna tecken.  
De här menykommandona väljer du genom att bara trycka på det understrukna tecknet.  
Dialogstyrning med tangentkombinationer  
I dialogrutor framhävs ett element i taget - som regel med en streckad kant.  
Man säger att det här elementet, som kan vara en kommandoknapp, ett alternativfält, en post i en listruta eller en kryssruta, är fokuserat.  
Om det fokuserade elementet är en kommandoknapp så utförs funktionen när du trycker på returtangenten, precis som om du hade klickat på knappen.  
Du markerar och avmarkerar en kryssruta genom att trycka på mellanslagstangenten.  
Om ett alternativfält är fokuserat växlar du till de andra alternativfälten i området med piltangenterna.  
Med Skift+Tabb hoppar du i motsatt riktning.  
Stäng en dialogruta med Esc om du inte vill göra några ändringar.  
En fokuserad kommandoknapp är inte bara omgiven av en streckad kant utan ofta också markerad med en något kraftigare skugga än de andra kommandoknapparna.  
Den kraftiga skuggan betyder följande:  
Om du stänger dialogrutan med hjälp av returtangenten är det detsamma som att trycka på den knapp som för tillfället är markerad med kraftigare skugga.  
Tangenter i kombination med musoperationer  
När du använder dra-och-släpp, markerar med musen samt klickar på objekt och namn startar du ytterligare funktioner med tangenterna Skift, Kommando Ctrl samt i enstaka fall Alternativ Alt.  
Tilläggsfunktionerna indikeras genom att muspekaren förändras när du samtidigt trycker på tangenter och använder dra-och-släpp.  
Tilläggstangenterna används bland annat till att utöka markeringen då du markerar filer, objekt, delar av text samt celler, rader och kolumner i tabeller.  
Funktionerna förklaras vid respektive beskrivning av de enskilda alternativen.  
Praktiska textinmatningsfält  
I alla textinmatningsfält och kombinationsfält där det går att göra inmatningar direkt har du tillgång till praktiska redigeringsmöjligheter.  
Prova det t.ex. i URL-fältet på funktionslisten:  
På en snabbmeny hittar du de mest använda kommandona.  
Med tangentkombinationen Skift + Kommando Ctrl +S öppnar du dialogrutan Infoga specialtecken.  
Med Kommando Ctrl +A markerar du hela textinnehållet.  
Med höger eller vänster piltangent tar du bort markeringen igen.  
När du dubbelklickar på ett ord markeras det.  
När du trippelklickar markeras hela innehållet.  
Med Kommando Ctrl +Delete raderar du från markörens position till slutet på det aktuella ordet.  
Håller du dessutom ner skifttangenten markerar du orden samtidigt.  
Med Insert växlar du mellan infogningsläge och överskrivningsläge.  
Du kan använda dra-och-släpp både innanför och mellan textfält.  
Med Kommando Ctrl +Z ångrar du ändringar steg för steg; texten har då samma innehåll som innan du gjorde den första ändringen.  
I %PRODUCTNAME finns AutoComplete-funktionen för en del text - och kombinationsfält.  
Om du t.ex. skriver c:\ i URL-fältet så visas den första filen eller katalogen på enheten C: (motsvarande för andra operativsystem) med hjälp av AutoComplete-funktionen.  
Nu kan du bläddra igenom alla andra filer och kataloger med hjälp av piltangenten Nedpil.  
Med Högerpil utökas visningen i URL-fältet till en eventuell underordnad katalog.  
En snabbare komplettering får du om du trycker på tangenten End så snart du har skrivit in en del av URL:en.  
När du har hittat ett program som du vill köra, eller ett dokument som du vill öppna, trycker du på returtangenten.  
Om du vill byta till en markerad katalog trycker du på returtangenten.  
Avbryta makron  
Om du vill avbryta ett aktivt makro trycker du på Skift + Kommando Ctrl +Q.  
Lista över allmänna tangentkombinationer i %PRODUCTNAME  
De tangentkombinationer som du kan använda i stället för menykommandon visas till höger om menytexterna på menyerna. (På Macintosh är inte alla tangenter som nämns tillgängliga för att styra dialogrutorna.)  
Tangentkombination  
Effekt  
Retur  
Motsvarar att du trycker på den fokuserade kommandoknappen i en dialogruta  
Esc  
Avbryter aktiviteten eller dialogrutan.  
I %PRODUCTNAME -hjälpen: hoppa tillbaka en nivå.  
Markören står i fältet URL på funktionslisten: markören placeras i dokumentet igen.  
Om en URL är markerad måste du trycka två gånger på tangenten.  
Blankstegstangent  
Växlar fokuserad kryssruta i en dialogruta  
Piltangenter  
Växlar aktivt kontrollfält i ett alternativområde i en dialogruta  
Tab  
Flyttar fokus till nästa område eller element i en dialogruta.  
Skift+Tab  
Flyttar fokus till föregående område eller till ett element i en dialogruta  
Alternativ Alt +Nedpil  
Öppnar listan för ett markerat kontrollfält i en dialogruta.  
Den här tangentkombinationen gäller både för kombinationsfält och för ikonknappar med popupmeny.  
Med Esc stänger du listan igen.  
Delete  
Raderar ett eller flera markerade objekt och placerar det / dem i papperskorgen  
Skift+Delete  
Raderar ett eller flera markerade objekt direkt (de placeras inte i papperskorgen)  
Backsteg (ovanför returtangenten)  
I en mappvy: gå upp en nivå (tillbaka)  
Kommando Ctrl +Tab  
Växlar till nästa öppnade dokument (utom i början av en överskrift: där infogas en tabulator)  
Skift + Kommando Ctrl +Tab  
Växlar till föregående öppnade dokument  
Kommando Ctrl +O  
Öppnar ett dokument  
Kommando Ctrl +S  
Sparar aktuellt dokument  
Kommando Ctrl +N  
Skapar nytt dokument  
Skift + Kommando Ctrl +N  
Öppnar dialogrutan Mallar och dokument  
Kommando Ctrl +P  
Skriver ut dokument  
Kommando Ctrl +Q  
Avslutar programmet  
Kommando Ctrl +X  
Klipper ut markerade element  
Kommando Ctrl +C  
Kopierar markerade element  
Kommando Ctrl +V  
Klistrar in från urklippet  
Kommando Ctrl +A  
Markerar allt  
Kommando Ctrl +Z  
Ångra  
Kommando Ctrl +G  
Öppnar dialogrutan Sök och ersätt.  
Kommando Ctrl +Skift+G  
Söker vidare efter det senast angivna sökordet.  
Ctrl+Skift+J  
Växlar mellan visning i helskärmsläge / normalläge  
Kommando Ctrl +Skift+R  
Uppdatering av dokumentfönstret  
Kommando Ctrl +K  
Det markerade området förses med attributet Kursiv.  
Om markören står i ett ord visas även det här ordet kursivt.  
Kommando Ctrl +F  
Det markerade området förses med attributet Fet.  
Om markören står i ett ord visas även det här ordet i fet stil.  
Kommando Ctrl +U  
Det markerade området förses med attributet Understrykning.  
Om markören står i ett ord blir även det här ordet understruket.  
Kommando Ctrl +Skift+O  
Sätter markören i fältet Ladda URL på funktionslisten.  
Alternativ Alt +O  
I dialogrutan för rättstavning överförs ordet som först var markerat som okänt / felaktigt (Original) till inmatningsraden (Ord).  
Några av de följande kombinationerna av funktionstangenter är inte tillgängliga för Mac.  
Tangentkombinationer med funktionstangenterna  
Tangentkombination  
Effekt  
F1  
Starta %PRODUCTNAME -hjälpen  
I %PRODUCTNAME -hjälpen: hopp till översiktssidan.  
Skift+F1  
Sammanhangsrelaterad hjälp  
Ctrl+F4 eller Alt+F4  
Stänger det aktuella dokumentet (stänger %PRODUCTNAME när det sista öppna dokumentet stängs)  
F6  
Sätter fokus i nästa delfönster (t.ex. dokument / datakällvy)  
Skift+F6  
Sätter fokus i föregående delfönster  
Skift+F10  
Öppnar snabbmenyn  
Tangentkombinationer inom plug-in-moduler  
I plug-in-moduler inom %PRODUCTNAME gäller följande tangentkombinationer:  
Tangentkombination  
Effekt  
F4  
Infogar hyperlänk  
F6  
Infogar OLE-objekt  
Support  
Sun Microsystems supportcentrum hjälper dig om du får problem med %PRODUCTNAME.  
Det finns en sammanfattning av alla supporttjänster som vi för närvarande erbjuder i en "Readme "-fil i %PRODUCTNAME -mappen.  
Besök vår hemsida på Internet, http: / /www.sun.com / staroffice, där du får mer information.  
På Sun Microsystems webbplats hittar du alltid aktuell information om Sun Microsystems och %PRODUCTNAME.  
Symboler i hjälpen  
Symboler i hjälpen  
De hänvisar till textavsnitt som innehåller mer information.  
Här följer en beskrivning av de enskilda symbolerna och deras betydelse.  
OBS!  
Den här symbolen hänvisar till ett textavsnitt som innehåller viktig information om data - och systemsäkerhet.  
Info!  
Det kan t.ex. beskriva ett annat sätt att göra samma sak.  
Tips!  
Den här symbolen visar att det finns ett tips om hur du kan arbeta ännu snabbare och effektivare med programmet.  
Hjälpfönstret i %PRODUCTNAME  
Observera att det här hjälpsystemet beskriver kommersiell programvara från Sun Microsystems, Inc.  
En del funktioner beskrivs visserligen här, men finns kanske inte med i den här %PRODUCTNAME -distributionen på grund av licensbegränsningar.  
Hjälpfönstret visar den valda sidan i hjälpen.  
Du kan visa och dölja ett navigationsområde.  
Symbollisten innehåller funktioner som är viktiga för hjälpsystemet:  
Aktivera / inaktivera navigationsområde  
Gå till föregående sida  
Gå till nästa sida  
Gå till startsidan i den aktuella hjälpen  
Skriva ut aktuell sida  
Lägg till bokmärke  
De här kommandona finns också på snabbmenyn (tryck på höger musknapp) i hjälpdokumentet.  
Om du vill kopiera från hjälpen till urklippet markerar du texten i hjälpen.  
Sedan väljer du Kopiera på snabbmenyn eller trycker på Kommando Ctrl +C.  
Med Tabb och Skift+Tabb växlar du mellan flikarna och hjälpdokumentet.  
Navigationsområde  
Navigationsområdet har flikarna Innehåll, Index, Sök och Bokmärken.  
Vid den övre kanten av området finns det en urvalslist där du kan välja hjälp till andra %PRODUCTNAME -moduler.  
Index och Sök refererar bara till den valda %PRODUCTNAME -modulen.  
Innehåll  
Under den här fliken finns en trädvy över huvudhjälpsidorna.  
Index  
Under den här fliken finns ett sorterat sakregister.  
Sök  
Under den här fliken kan du göra en textsökning i hela hjälpinnehållet i den valda %PRODUCTNAME -modulen.  
Bokmärke  
Den här fliken innehåller de bokmärken som du har definierat.  
Här kan du redigera och radera definierade bokmärken eller byta till motsvarande sida.  
Help Agent, tipshjälp och aktiv hjälp  
De här funktionerna kan du använda i programmet utan att behöva aktivera hjälpfönstret.  
Välj på menyn Hjälp.  
Help Agent  
Help Agent öppnas automatiskt i vissa situationer.  
Om du klickar på fönstret får du hjälp till den aktuella situationen.  
Tipshjälpen  
Håll markören över en kommandoknapp så visar tipshjälpen namnet på kommandoknappen.  
Dessutom visar tipshjälpen annan information på många ställen, t.ex. kapitelnamn när du rullar genom ett långt dokument.  
Den aktiva hjälpen  
Om du vill få en kort beskrivning av en funktion hos en kommandoknapp, ett inmatningsfält eller ett menykommando väljer du den aktiva hjälpen.  
Du aktiverar även den här funktionen via Skift+F1.  
Index - nyckelordssökning i hjälpen  
Ange ett ord i indexlistan eller dubbelklicka på en post.  
Här visas en lista i två nivåer med indexord för det valda programområdet.  
Klicka här för att visa det valda ämnet.  
Här kan du söka efter ett specifikt ämne.  
I det undre fönstret ser du en alfabetiskt ordnad lista över alla indexposter.  
I det övre inmatningsfältet Sökord kan du söka efter ett specifikt ord i indexlistan.  
Om markören är placerad i Indexlistan hoppar du direkt till nästa passande post när du matar in ett sökord.  
Om du matar in ett sökord i inmatningsfältet Sökord hoppar du till motsvarande post i indexlistan så snart ett ord hittas som motsvarar sökordet.  
Hjälpindex och textsökning gäller alltid det område som har valts senast i %PRODUCTNAME.  
Om du inte får något sökresultat bör du först kontrollera om du har valt rätt hjälpområde.  
Söka - textsökningen  
Mata in sökordet här.  
Sökningen tar inte hänsyn till skrivsätt med stor eller liten bokstav.  
Klicka här när du vill starta textsökningen efter det angivna sökordet.  
Här visas rubrikerna på de hittade sidorna som resultat av din textsökning, sorterat efter relevans med de bästa träffarna i början av listan.  
Om du vill titta på en sida dubbelklickar du på posten.  
Markera den här rutan om du vill göra en exakt sökning efter det angivna sökordet.  
Delar av ord hittas inte.  
Markera den här rutan om du bara vill söka i dokumentrubriker.  
Klicka här om du vill se den markerade posten i träfflistan.  
Textsökningsfunktionen i %PRODUCTNAME -hjälpen gör att du kan hitta hjälpdokument som innehåller olika kombinationer av sökord.  
Mata in ett eller flera ord i inmatningsfältet Sökord.  
Inmatningsfältet Sökord kommer ihåg de senast inmatade sökorden.  
Du kan välja dem igen från listan om du vill upprepa sökningen.  
När sökningen är avslutad visas rubrikerna på de hittade dokumenten i listan, sorterade i fallande ordning efter relevans, d.v.s. med de bästa träffarna längst upp.  
Du laddar ett hjälpdokument genom att dubbelklicka på en post eller genom att markera en post och klicka på Visa.  
Med hjälp av Sök bara i rubriker kan du begränsa sökningen till dokumentrubriker.  
Kryssrutan Bara hela ord gör att du kan göra en exakt sökning.  
Om den här rutan är markerad hittas inga delar av ord.  
Markera inte den här rutan om det angivna sökordet även ska hittas som del av ett längre ord.  
Du kan använda en valfri kombination av sökord, åtskiljda med mellanslag.  
Sökningen är inte versalkänslig.  
Hjälpindex och textsökning gäller alltid det program som har valts senast.  
Om din sökning inte ger något resultat bör du först kontrollera att du har valt rätt hjälpområde.  
Administrera bokmärken  
Här kan du ange ett nytt namn för bokmärket vid behov.  
Med ikonen Lägg till bokmärke sätter du ett bokmärke på sidan som visas i hjälpen.  
Bokmärkena visas under fliken Bokmärken.  
Om du dubbelklickar på ett bokmärke eller trycker på returtangenten öppnas den tilldelade sidan i hjälpen.  
Om du klickar med höger musknapp öppnas snabbmenyn.  
Du raderar det valda bokmärket med Delete-tangenten utan säkerhetskontroll.  
I snabbmenyn till ett bokmärke finns det följande kommandon:  
Visa - visar det markerade ämnet i hjälpen.  
Byt namn - öppnar en dialogruta där du matar in ett annat namn för bokmärket.  
Radera - raderar det markerade bokmärket.  
Innehåll - huvudämnena i hjälpen  
Här ser du huvudämnena i hjälpen i en struktur som liknar mapparna i en filhanterare.  
Dubbelklicka på en stängd mappsymbol om du vill öppna mappen och visa de underordnade mapparna och hjälpsidorna som finns i den.  
Dubbelklicka på en öppen mappsymbol om du vill stänga mappen och dölja de underordnade mapparna och hjälpsidorna som finns i den.  
Dubbelklicka på en dokumentsymbol om du vill öppna motsvarande hjälpsida.  
Med piltangenterna i kombination med returtangenten kan du öppna och stänga poster och öppna dokument.  
Hjälpsidan hittades inte.  
Tyvär gick det inte att hitta hjälpsidan som du har valt.  
Följande data kan vara till hjälp när felet ska identifieras:  
Hjälp-ID:  
<help:error-id xmlns:help=" http: / /openoffice.org / 2000 / help "/ >  
Hjälpmodul:  
<help:error-module xmlns:help=" http: / /openoffice.org / 2000 / help "/ >  
Hjälpsökväg:  
<help:error-path xmlns:help=" http: / /openoffice.org / 2000 / help "/ >  
Det här felmeddelandet kan ha följande orsaker:  
Hjälpmodulen är inte installerad.  
Vid installationen kan du välja vilka hjälpmoduler som ska installeras.  
Om du inte har installerat alla hjälpmoduler eller program har hjälpsystemet inte tillgång till motsvarande fil.  
Så ändrar du en existerande installation.  
Databasen för hjälptexten är skadad.  
Filerna för hjälptexterna administreras via en databas.  
Den kan ha blivit skadad antingen på grund av en skadad installation eller egna ändringar.  
Så här reparerar du en skadad installation.  
Klicka på Tillbaka om du vill gå tillbaka till den föregående sidan.  
Skapa en hemsida  
Här ser du hur du skapar en egen hemsida för Internet och ger den en intressant grafisk utformning med olika hjälpmedel i %PRODUCTNAME.  
Till slut måste du lägga upp hemsidan hos en Internet-leverantör och registrera den hos olika sökmotorer.  
Så här gör du i ordning en hemsida på Internet:  
Skapa sidan (sidorna) i %PRODUCTNAME.  
Utforma eller sök efter de grafiska objekt som du vill ha med på sidan och arkivera alla som filer i en katalog.  
Det är bäst att använda katalogen där dina HTML-textfiler finns eller en underordnad katalog till den.  
Du bör även spara använda grafiska objekt från Gallery som egna filer.  
Infoga de grafiska elementen som länkar i %PRODUCTNAME -textdokumenten.  
Kontrollera hur sidorna ser ut och fungerar med olika webbläsare.  
Ladda sidorna till utrymmet för din hemsida hos din Internet-leverantör.  
Du kan använda den som utgångspunkt för din egen sida.  
Så här utformar du en egen hemsida med %PRODUCTNAME.  
Den hjälper dig interaktivt; de enskilda stegen förklaras i beskrivningen av Arkiv - AutoPilot.  
Ge HTML-sidan en rubrik!  
Den visas på titellisten i webbläsare när en besökare tittar på din sida och används även som bokmärke.  
Rubriken skriver du in i dialogrutan Arkiv - Egenskaper - Beskrivning i fältet Rubrik.  
Spara den här sidan som HTML-fil i en katalog som du har reserverat för filer som hör till hemsidan.  
Katalogen kan t.ex. heta "C: \hemsida".  
Här samlar du alla filer som hör till din hemsida och kan senare överföra alla till din Internet-leverantör samtidigt.  
Mata in namnet "Start.htm" eller "Index.htm ".  
Fråga din Internet-leverantör om den första sidan (startsidan) på din hemsida måste ha ett särskilt namn för att den ska laddas automatiskt, utan att sidan behöver anges.  
Kontrollera nu att URL:erna på dina sidor sparas i filsystemet med relativa sökvägar.  
Det är viktigt för att länkarna till andra element på hemsidan ska kunna fungera i varje katalog och på varje enhet.  
Markera rutan i filsystem i området Spara URL:er relativt under Verktyg - Alternativ - Ladda / spara - Allmänt.  
Hemsidans katalogstruktur  
För att du ska kunna infoga grafik utan problem på din HTML-sida på leverantörens server bör du tänka på följande:  
Skapa en mapp för din hemsida på hårddisken.  
Kalla den t.ex. för "hemsida".  
Det är alltså här som du sparar din HTML-startfil som vanligen bör heta "index.htm".  
Kalla t.ex. den underordnade katalogen för "grafik". (Det är bra att genomgående skriva alla fil - och mappnamn med små bokstäver eftersom det finns servrar som hanterar filer och mappar olika beroende på om de är skrivna med stora eller små bokstäver.)  
Skapa även en underordnad katalog med namnet "grafik" i området för din hemsida på leverantörens server.  
Länka bara till grafik som ligger i den underordnade katalogen "grafik" på dina HTML-sidor.  
Det gör du genom att integrera relativa länkar av typen <IMG SRC=" grafik / bild1.gif ">.  
Detta förutsätter att all grafik har infogats som länkar och att du redan har konverterat all grafik till GIF - eller JPG-format. %PRODUCTNAME kan visserligen också omvandla inbäddad grafik till GIF-filer automatiskt och infoga motsvarande taggar på HTML-sidan.  
Men då har du ingen kontroll över filnamnen och för grafik som du har lagt in på flera ställen skapas det också flera filer.  
Testa din hemsida lokalt.  
Ladda även all grafik från den lokala mappen "grafik" till mappen med samma namn hos leverantören.  
Integrera grafik på hemsidan  
När du arbetar med din hemsida bör du växla till onlinelayout-läge, om du inte har börjat direkt med ett %PRODUCTNAME Writer / Web-dokument.  
Då kan du bara utföra kommandon som leder till sidelement som är tillåtna i HTML-läge.  
Du växlar till onlinelayout på Visa -menyn.  
Grafik som ska användas på Internet måste vara i GIF - eller JPG - (eller PNG -) format.  
Integrerad grafik i andra format skulle %PRODUCTNAME automatiskt omvandla till JPG-format när den exporteras som HTML-dokument.  
För att du ska få en välstrukturerad och lättskött hemsida är det i varje fall bättre om du själv gör konverteringen till GIF eller JPG.  
Öppna %PRODUCTNAME och ladda ett grafikobjekt.  
Spara grafikobjektet med Arkiv - Spara som i filformatet GIF eller JPG, helst i en underordnad katalog till C:\hemsida (se ovan),.  
Stäng %PRODUCTNAME.  
Sätt markören på det ställe på hemsidan där du vill infoga ett grafikobjekt.  
Välj JPG-grafiken från hemsideskatalogen under Infoga - Grafik - Från fil och markera fältet Länka.  
Klicka på kommandoknappen Öppna så infogas grafikobjektet.  
Annars kan du få oönskade effekter (trappstegseffekt vid förstoring, problem med tunna linjer vid förminskning o.s.v.).  
Ändra bakgrund för hemsida  
Klicka på ett ledigt utrymme på sidan så att bilden inte längre är markerad.  
Öppna dialogrutan Format - Sida och klicka på fliken Bakgrund.  
I listrutan som väljer du Färg.  
Välj en annan bakgrundsfärg och klicka på OK.  
Om du skulle välja Grafik i listrutan kan du lägga in ett bakgrundsgrafikobjekt - det kan du prova nästa gång.  
Sedan kan du välja om bakgrundsgrafikobjektet ska placeras centrerat, vid en kant eller upprepade gånger sida vid sida så att hela bakgrunden täcks.  
Överföra filerna för hemsidan till Internet-leverantören  
När hemsidan ser ut precis som du vill ha den, kan du överföra alla filer från hemsideskatalogen till utrymmet för din hemsida hos Internet-leverantören.  
Detaljerade anvisningar får du av leverantören.  
Skapa en enkel hemsida  
Om du snabbt vill lägga upp en hemsida med grafik på Internet kan du göra det utan allt för mycket förarbete:  
Öppna en ny, tom sida för hemsidan (med Arkiv - Nytt - HTML-dokument).  
Lägg in bilder som du vill (som länkar eller direkt inbäddade objekt, via dialogrutan Infoga - Grafik eller genom att dra dem från Gallery och släppa dem i HTML-dokumentet).  
Spara dokumentet lokalt.  
Men det behöver du inte bekymra dig om i det här läget.  
Öppna dialogrutan Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet och kontrollera att rutan Kopiera lokal grafik till Internet är markerad.  
Anslut till Internet.  
Spara sidan med dialogrutan Arkiv - Spara som...  
Ange hemsidans fullständiga URL hos leverantören i fältet Filnamn, t.ex. enligt mönstret http: / /hemsidor.leverantör.com / mittnamn / index.htm.  
Nu konverterar %PRODUCTNAME automatiskt all länkad och inbäddad grafik på sidan till GIF-format.  
Grafikobjekten får nya, entydiga namn.  
I HTML-dokumentet skapas länkar till grafikobjekten enligt mönstret <IMG SRC=" abc123.gif ">, alltså med relativ sökväg.  
HTML-sidan och all grafik överförs sedan till den angivna katalogen.  
HTML-mallen i %PRODUCTNAME  
Om du vill skapa en ny sida för Internet öppnar du ett nytt HTML-dokument under Arkiv - Nytt.  
När du skriver Internet-sidor är det även till god hjälp att använda onlinelayout-läget, som du kan aktivera på menyn Visa.  
I onlinelayout-läget har du bara tillgång till de menyer och dialogrutor i %PRODUCTNAME som gäller för HTML-sidor.  
Skapa en ny sida för Internet  
Växla först till Onlinelayout-läge genom att markera det alternativet på Visa -menyn eller påbörja ett nytt HTML-dokument. %PRODUCTNAME använder då internt formatmallen html.vor som finns i mappen {installpath} / share / template / swedish / internal.  
På den nya sidan kan Du skriva in text, infoga objekt osv precis som på "normala" sidor.  
Använd de särskilda stycke - och teckenformatmallar som redan finns i HTML-mallen.  
Vid intern export till HTML försöker %PRODUCTNAME dessutom bibehålla originaldokumentet intakt så långt möjligt inom ramen för HTML-formatet.  
Om du vill göra om ett %PRODUCTNAME -dokument till en HTML-sida sparar du sidan i filformatet Webbsida.  
Ge filen ett namn som slutar med filnamnstillägget .HTM eller .HTML.  
Sidformatmall HTML (normal)  
I den här sidformatmallen används inga marginaler för sidorna och sidorna kan göras nästan hur långa som helst utan störande sidbrytningar.  
Styckeformatmallar för HTML-sidor  
De särskilda styckeformatmallarna för HTML-sidor har följande egenskaper:  
Styckeformatmall  
Betydelse  
BLOCKQUOTE  
Citat kan formateras som BLOCKQUOTE.  
Texten visas då t ex med indrag och i kursiv stil.  
DD 1-3, DT 1-3  
Ordlistor kan struktureras med hjälp av DT - och DD-format.  
Första nivån definieras som första ordlistetemat med DT1 och tillhörande text definieras med DD1.  
Rubriken på första undernivån får formatet DT2 och texten får formatet DD2.  
Tredje nivån får på motsvarande sätt formatet DT3 och DD3.  
Indragen görs så att DT1 står längst till vänster, DD1 dras in ett steg, DT2 dras in till samma nivå som DD1 osv.  
HR  
En horisontell linje infogas över hela sidans bredd.  
PRE  
Texten formateras som "förformaterad text" i teckensnittet Courier med fasta breddsteg.  
Eftersom alla blanksteg även visas i HTML-text, är det här formatet lämplig för programförteckningar etc som dras in med blanksteg.  
Teckenformatmallar för HTML-sidor  
Även de särskilda teckenformatmallarna för HTML-sidor (Du kan givetvis även använda andra formatmallar) anges med versaler.  
Följande teckenformatmallar finns:  
Teckenformatmall  
Betydelse  
Internet-länk  
Tecknen formateras i blått med understrykning  
använd Internet-länk  
Tecknen formateras i rött med understrykning  
ABBREV  
logisk effekt för förkortningar  
ACRONYM  
logisk effekt för akronymer (ord som består av begynnelsebokstäverna i andra ord)  
AU  
logisk effekt för författarnamn  
BLINK  
logisk effekt för blinkande text  
CITE  
logisk effekt för citat (t.ex. kursiv stil)  
CODE  
logisk effekt för källkod (t.ex. Courier)  
DEL  
logisk effekt för raderad text (ändringsmarkering)  
DFN  
logisk effekt för en definition  
EM  
logisk effekt för framhävning (t.ex. kursiv stil)  
INS  
logisk effekt för infogad text (ändringsmarkering)  
KBD  
logisk effekt för skärmtecken (t.ex. Courier)  
LANG  
logisk effekt för främmande språk  
PERSON  
logisk effekt för personnamn  
Q  
logisk effekt korta citat  
SAMP  
logisk effekt för exempel (t.ex. Courier)  
STRONG  
logisk effekt för viktig text (t.ex. fet stil)  
TT  
logisk effekt för teckensnitt med fasta breddsteg (t.ex. Courier)  
VAR  
logisk effekt för variabel (t.ex. kursiv stil)  
Flera av dessa formateringar inkluderas med HTML-taggar vid export till HTML-format, men visas som normal text av många webbläsare.  
Formateringar som omvandlas till HTML  
%PRODUCTNAME kan t ex skapa en lämplig HTML-kod med utgångspunkt från ett %PRODUCTNAME -textdokument.  
Uppräkningar exporteras t ex i ett textdokument som HTML-taggar som kan visas som en uppräkning eller lista i webbläsaren.  
I följande lista redovisas en del av dessa formateringar:  
Formatering i ett %PRODUCTNAME -dokument  
Typ av HTML-tagg som skapas  
(Huvudet skapas automatiskt)  
<head>  
Titel i dialogrutan Dokumentegenskaper  
<titel>  
Styckeformatmallarna Överskrift 1 till x  
<H1> till <Hx>  
Styckeformatmall Avsändare  
<address>  
Tabell i textdokument  
<table ...>  
Attributet fet  
<b>  
Attributet kursiv  
<i>  
Attributet understrykning  
<u>  
Punktlistor (punktuppställning)  
<ul> som inledning, <li> för varje listelement  
Numreringar  
<ol> som inledning, <li> för varje listelement  
Index (nedsänkning)  
<sub>  
Exponent (upphöjning)  
<super>  
infogad anteckning  
<!- - blir en kommentar -->  
infogat område  
<div ID=" områdesnamn ">.....< / div>  
AutoKorrigering har aktiverats  
TVå versaler i ordets början korrigerades.  
Skrivfel som "ORd" korrigeras till "Ord "av AutoKorrigering.  
AutoKorrigering har aktiverats  
Börja varje mening med stor bokstav.  
Din text har korrigerats av AutoKorrigering: varje ord efter slutet på en mening (representerat av t.ex. punkt, utropstecken, frågetecken) börjar med stor bokstav.  
AutoKorrigering har aktiverats  
Två stora bokstäver i början av ett ord och i början av en mening korrigerades till en versal  
Din text korrigerades av AutoKorrigering: två stora bokstäver i början av ordet samt i början av meningen ersätts av en versal  
AutoKorrigering har aktiverats  
AutoKorrigering (en ersättning) utfördes  
AutoKorrigering gjorde en ersättning  
AutoKorrigering har aktiverats  
AutoKorrigering (ersättning) utfördes, meningen inleds nu med stor bokstav  
AutoKorrigering ersatte en bokstav så att meningen börjar med stor bokstav  
AutoKorrigering har aktiverats  
Dubbla citattecken har ersatts  
Din text korrigerades av AutoKorrigering: dubbla citattecken har ersatts av typografiska citattecken.  
AutoKorrigering har aktiverats  
Enkla citattecken har ersatts  
Din text har korrigerats av AutoKorrigering: enkla citattecken har ersatts av typografiska citattecken.  
AutoKorrigering har aktiverats  
En URL identifierades och försågs med hyperlänk-attribut  
Din text korrigerades av AutoKorrigering: en teckensträng identifierades som URL och visas nu som hyperlänk.  
AutoKorrigering har aktiverats  
Dubbla blanksteg ignorerades  
Din text korrigerades av AutoKorrigering: flera mellanslag efter varandra har sammanfattats till ett enda mellanslag.  
AutoKorrigering har aktiverats  
Fet eller understruken text identifierades och tilldelades  
Din text korrigerades av AutoKorrigering: textattributen fet och / eller understruken har tilldelats automatiskt.  
AutoKorrigering har aktiverats  
1 / 2... ersattes med ½...  
Din text har korrigerats av AutoKorrigering: en teckenkombination som motsvaras av ett enda tecken i teckenuppsättningen, t.ex. 1 / 2, har ersatts av respektive tecken.  
AutoKorrigering har aktiverats  
Tankstreck ersattes  
Din text korrigerades av AutoKorrigering: ett minustecken har ersatts av ett tankstreck.  
AutoKorrigering har aktiverats  
1st... ersattes med 1^st...  
Din text korrigerades av AutoKorrigering: de engelska ordningstalen, där slutet på talet placeras högre upp, har använts.  
AutoPilot  
Med hjälp av AutoPiloten utformar du egna dokumentmallar för affärsbrev och privata brev, fax, PM, presentationer och mycket annat.  
Brev...  
Fax...  
Agenda...  
PM...  
Presentation...  
Webbsida...  
Formulär  
Dokumentkonverterare  
Eurokonverterare...  
%PRODUCTNAME 5.2 databasimport  
Om du får ett felmeddelande om att "rättigheter saknas" när du försöker utföra en AutoPilot så har du troligen angett att Basic-makron aldrig ska utföras under Verktyg - Alternativ - %PRODUCTNAME - Säkerhet.  
Ändra inställningen från utför aldrig till utför alltid eller enligt lista.  
AutoPilot Brev  
Den kan användas som mall både för privata brev och affärskorrespondens.  
%PRODUCTNAME har en mönstermall för privata brev och affärskorrespondens, som du kan anpassa efter din personliga smak med hjälp av AutoPiloten.  
AutoPiloten leder dig steg för steg genom de olika layoutelementen i dokumentmallen och ger dig möjlighet att välja olika alternativ i varje steg.  
Den förminskade förhandsvisningen i dialogrutan ger dig ett första intryck av vilken effekt de aktuella inställningarna har.  
I dialogrutan kan du när som helst ångra ett val eller hoppa över enskilda eller alla steg.  
Om du hoppar över ett eller flera steg använder AutoPiloten de aktuella standardinställningarna.  
På sidan 5 i dialogrutan kan du göra inställningar för affärsbrev.  
De här inställningarna används normalt inte för privata brev, som t.ex. en ärendemening.  
För privata brev står dessutom mottagaren bara på kuvertet, inte på brevets förstasida.  
Därför saknas sidorna 4 och 5 i dialogrutan om du väljer alternativet Privat brev här.  
AutoPilot Brev - sida 2  
AutoPilot Brev - sida 6  
AutoPilot Brev - sida 8  
<< Tillbaka  
I dialogrutan kan du titta på urvalet i steget innan.  
De aktuella inställningarna finns kvar.  
Den här kommandoknappen är bara tillgänglig fr.o.m. det andra redigeringssteget.  
Nästa >>  
När du klickar på den här kommandoknappen använder AutoPiloten de aktuella inställningarna i dialogrutan och fortsätter till nästa steg.  
Om du har kommit till det sista steget i dialogrutan går det inte längre att välja den här kommandoknappen.  
Färdigställ  
AutoPiloten skapar en ny dokumentmall enligt dina inställningar och sparar den på hårddisken. %PRODUCTNAME skapar ett nytt dokument med namnet "namnlösX" (X står för ett löpnummer) som baserar på den nya dokumentmallen och visar det i arbetsområdet.  
%PRODUCTNAME sparar de aktuella inställningarna i AutoPiloten för den använda malltypen och använder dem som förinställningar nästa gång du startar AutoPiloten.  
AutoPilot Brev - sida 1  
På första sidan anger du om du vill skriva ett privat brev eller ett affärsbrev.  
Ditt val styr vilka alternativ som är tillgängliga på de följande sidorna.  
Vilken typ av brevmall vill Du skapa?  
Välj här om du vill skapa en mall för ett privat brev eller ett affärsbrev.  
Affärsbrev  
Välj det här alternativet, om du t.ex. behöver en ärenderad.  
Privat brev  
För ett privat brev skapas en mindre formell mall.  
Vilken stil vill Du använda?  
Här väljer du en av följande stilar för din brevmall:  
Modern Klassisk och Elegant.  
Du kan även titta på mallen på prov så att du ser hur den ter sig.  
Modern  
Här används främst teckensnitt utan seriffer.  
Klassisk  
Här används främst icke-proportionella teckensnitt.  
Elegant  
Här används främst antikvateckensnitt (med seriffer).  
Gå vidare till AutoPilot Brev - sida 2  
AutoPilot Brev / Fax - sida 2  
I det här området väljer du en logotyp för din mall.  
Beroende på vilken logotyp du väljer ändras de tillgängliga alternativen på den här sidan.  
Vilken typ av logotyp vill Du ha på brevet / faxet?  
I det här området väljer du en logotyp.  
Beroende på vilken slags logotyp du väljer ändras de tillgängliga alternativen på den här sidan.  
Ingen logotyp  
Markera det här alternativfältet om du inte vill ha någon logotyp på brevet / faxet.  
Ändringen visas symboliskt i förhandsvisningsfältet.  
Grafik  
Markera det här fältet om du vill ha ett grafikobjekt som logotyp.  
I området Grafikfilnamn kan du sedan välja en grafikfil.  
Text  
Markera det här fältet om du vill använda en text som logotyp.  
Storlek och teckensnitt kan du ändra senare.  
Grafikfilnamn  
Det här alternativet är bara synligt om du valt ett grafikobjekt som logotyp.  
Namnet på den valda grafikfilen visas; du kan välja en ny fil med kommandoknappen Grafikurval.  
Grafikurval...  
Med den här kommandoknappen öppnar du dialogrutan Välj logotypgrafik.  
Logotyptext  
Om du har valt en text som logotyp visas det flerradiga textfältet Logotyptext.  
Här matar du in den text som ska visas som logotyp i brevet.  
Storlek  
I området Storlek väljer du exakt numerisk storlek för logotypen i två rotationsfält, oavsett om logotypen utgörs av text eller grafik.  
Bredd  
Ställ in logotypens bredd här.  
Höjd  
Ställ in logotypens höjd här.  
Position  
Du kan finjustera positionen med rotationsfälten:  
Till vänster  
Med den här kommandoknappen placerar Du logotypen till vänster.  
Centrerat  
Med den här kommandoknappen placerar Du logotypen i mitten.  
Till höger  
Med den här kommandoknappen placerar Du logotypen till höger.  
Från vänster / höger  
Här kan du ställa in avståndet från logotypen till vänster eller höger sidmarginal.  
Uppifrån  
Här kan du ställa in avståndet från logotypen till den övre sidmarginalen.  
Gå vidare till AutoPilot Brev - sida 3  
Gå vidare till AutoPilot Fax - sida 3  
AutoPilot Brev - sidan 3  
På den här sidan bestämmer du hur brevet ska se ut och vad som ska stå i avsändaruppgifterna.  
Ange nu avsändaren:  
I det här textfältet anger du avsändaruppgifterna.  
I denna form kommer de sedan att visas som redigerbar text i alla brev som du skriver med hjälp av den här brevmallen.  
Du kan därför trycka på returtangenten vid varje radslut i det här fältet utan att dialogrutan stängs.  
Lägg märke till att det första tecknet i adressfönstret måste vara ">".  
Alla rader som börjar på det sättet upprepas i mottagarfältet, såvida du tillåter det generellt (se nästa fält).  
Uppdatera adress från användardata  
Genom att klicka på den här symbolen ersätter du texten i avsändarfältet med en standardinställning för avsändare, som baseras på användardata.  
Upprepa i mottagarfält?  
Här kan du bestämma om avsändaren ska anges i liten stil ovanför mottagaren, så att den går att läsa i ett fönsterkuvert.  
Ja  
Om du gör en markering här, visas de avsändarrader som börjar med ">" i mottagarfältet.  
Nej  
Om du gör en markering här, visas avsändaren inte i mottagarfältet.  
Position och storlek  
Med hjälp av alternativfälten, som innehåller en liten förhandsvisning av avsändarens position, kan du på ett ungefär ange positionen för avsändarfältet.  
Sedan kan du ställa in exakt med rotationsfälten.  
Uppe till vänster  
Här hamnar avsändaren uppe till vänster på sidan.  
Uppe till höger  
Här hamnar avsändaren uppe till höger på sidan.  
Nere till vänster  
Här hamnar avsändaren nere till vänster på sidan.  
Nere till höger  
Här hamnar avsändarfältet nere till höger på sidan.  
Till höger bredvid mottagaren  
Här hamnar avsändaren till höger om mottagaren på sidan.  
Från vänster / höger  
Här definierar Du avståndet mellan avsändarfältet och den vänstra eller högra sidmarginalen.  
Uppifrån / nerifrån  
Här definierar du avståndet mellan avsändarfältet och den undre sidmarginalen.  
Bredd  
Här ställer du in avsändarfältets bredd.  
Höjd  
Här ställer du in avsändarfältets höjd.  
Gå vidare till AutoPilot Brev - sidan 4  
AutoPilot Brev - sida 4  
På den här sidan kan du definiera databastypen och databasfält för hälsningsfrasen.  
Databas  
Här väljer du databasen som innehåller poster för mottagaruppgifterna.  
Databas  
Här väljer du den tabell där mottagaruppgifterna ska hämtas i den aktuella databasen.  
Posterna i den här listrutan ändras beroende på urvalet i den vänstra listrutan Databas.  
Adress  
Här sammanställer Du uppgifterna om mottagaren.  
Mottagarens adress kan Du antingen skriva in direkt - sedan står den alltid så i mallen - eller så kan Du ange databasfält som används som platshållare för innehåll från databasen.  
Fördelen med detta är att Du direkt kan använda mallen till att skriva ut standardbrev.  
Databasfält  
Här väljer Du genom att klicka på ett fält som Du vill överföra till mottagarfältet.  
Vänsterpil  
Klicka på den här pilen om det markerade databasfältet vid markörens aktuella position ska överföras till fältet Adress.  
Styckebrytning  
Klicka här om Du vill infoga en styckebrytning vid markörens aktuella position i adressfältet.  
Du kan också trycka på Retur i stället.  
Hälsningsfras  
I fälten till hälsningsfrasen kan Du ange ett tilltal som ska infogas framför brevets textområde.  
I listrutan kan Du välja ett av databasens fält, vars innehåll ska överföras till raden med hälsningsfrasen (t.ex. förnamn).  
Tilltalet kan du också bara definiera via listrutan, om databasen t.ex. innehåller ett fält för Tilltal.  
Gå vidare till AutoPilot Brev - sida 5  
AutoPilot Brev - sida 5  
På den här sidan definierar du vilka layoutelement ditt dokumentet ska innehålla.  
Markera rutan bredvid det element som du vill använda.  
1.  
Er referens  
Markera den här rutan om du vill använda standardelementet Er referens i din text.  
Er referens  
Du kan redigera texten vid behov, eller överta standardelementet i ditt brev.  
2.  
Vår referens  
Markera den här rutan om du vill använda standardelementet Vår referens i din text.  
Vår referens  
Överta standardtexten eller redigera den enligt dina önskemål.  
3.  
Ert brev daterat  
Markera den här rutan om du vill använda standardelementet Ert brev daterat i din text.  
Ert brev daterat  
Överta standardtexten eller redigera den.  
4.  
Vårt brev daterat  
Markera den här rutan om du vill använda standardelementet Vårt brev daterat i din text.  
Vårt brev daterat  
Använd standardtexten eller redigera den enligt dina önskemål.  
Datum  
Markera den här rutan om du vill infoga dagens datum som fältfunktion i din brevmall.  
Datum  
Här väljer du datumformat.  
Ärenderad  
Markera den här rutan om du vill infoga en ärenderad.  
Ärenderad  
Här skriver du texten för ärenderaden.  
Kopia till  
Markera den här rutan om du vill använda texten Kopia till i din brevmall.  
Bilaga / or  
Markera den här rutan om du vill använda texten Bilaga / or i din brevmall.  
Sidnummer  
Markera den här rutan om du vill ha sidnummer i din brevmall.  
I de följande fälten kan du sedan bestämma hur sidnumret ska anges.  
"Sida"  
Här skriver du den text som ska skrivas ut framför sidnumret. "Sida" är fördefinierat.  
Listrutan Sidnummer  
I den här listrutan väljer du den stil med vilken sidorna ska numreras.  
Totalt antal sidor  
Markera den här rutan om även det totala sidantalet i brevet ska nämnas i området med sidnummer.  
Textfältet Totalt antal sidor "av"  
I förinställningen visas sidantalet enligt mönstret Sida x av y.  
Texten av kan du ändra i det här textfältet om du vill, t.ex. ersätta den med /.  
Gå vidare till AutoPilot Brev - sida 6  
AutoPilot Brev / Fax - sida 6  
På den här sidan definierar du utseendet för sidfoten och bredden på sidmarginalerna.  
Sidfot  
I det här området kan du mata in en sidfot som infogas på varje sida i ditt brev / fax.  
Sidfot på  
Markera det här fältet för att infoga en sidfot.  
Skiljelinje för text  
Markera den här rutan om du vill infoga en skiljelinje mellan text och sidfot.  
Nerifrån (bara för brev)  
Här anger du avståndet mellan sidfoten och den undre sidmarginalen.  
Till text (bara för brev)  
Här anger du avståndet mellan sidfot och text.  
Sidfot  
I det här flerradiga textfältet matar du in text för sidfoten.  
Sidmarginaler  
I förhandsvisningen kan du se effekten av de här inställningarna.  
Från vänster  
Här definierar du den vänstra sidmarginalen.  
Från höger  
Här definierar du den högra sidmarginalen.  
Gå vidare till AutoPilot Brev - sida 7  
Gå vidare till AutoPilot Fax - sida 7  
AutoPilot Brev - sidan 7  
Här definierar du utseendet på de efterföljande sidorna.  
Sidhuvud  
I det här området definierar du layouten för ditt sidhuvud.  
Det kan innehålla logotypen och avsändaren.  
Uppifrån  
Här anger du avståndet mellan sidhuvudet och den övre kanten på sidan.  
Tänk på det icke utskrivbara området (som bestäms av skrivarens egenskaper).  
Till text  
Här anger du sidhuvudets avstånd från den följande texten.  
Logotyp  
Här väljer du om och var logotypen ska upprepas.  
Du kan ställa in en annan storlek på logotypen för de följande sidorna än för den första sidan.  
Bredd  
Här ställer du in logotypens bredd.  
Höjd  
Här ställer du in logotypens höjd.  
Avsändare  
Du kan ställa in en annan storlek på avsändarfältet för de följande sidorna än för den första sidan.  
Bredd  
Här ställer du in avsändarfältets bredd.  
Höjd  
Här ställer du in avsändarfältets höjd.  
Sidfot  
I det här området anger du om och var sidfoten ska upprepas på de följande sidorna.  
Visa sidfot  
Klicka i den här rutan när du vill visa resp. dölja sidfoten.  
Nerifrån  
Här anger du avståndet mellan sidfoten och den nedre kanten på sidan.  
Ta hänsyn till det icke utskrivbara området (som bestäms av skrivarens egenskaper).  
Till text  
Här anger du avståndet mellan sidfoten och texten som ligger ovanför.  
Gå vidare till AutoPilot Brev - sidan 8  
AutoPilot Brev - sida 8 / Fax - sida 7 / PM - sida 4 / Agenda - sida 5  
På den här sidan definierar du var och med vilket namn dokumentet och dokumentmallen ska arkiveras.  
Dokumentinformation  
Här definierar du vilka uppgifter som ska finnas i dokumentegenskaperna (menyn Arkiv - Egenskaper) för dokument som skapas med den här mallen.  
Det går bara att välja inställningarna i det här området om du skapar en mall för affärsbrev, inte för privata brev.  
För kopplade utskrifter kan du även ange att innehållet i ett databasfält ska infogas som dokumentinfomation för varje enskilt dokument.  
Rubrik  
Här kan du välja det datafält, vars innehåll ska infogas som rubrik i dialogrutan Egenskaper  
Ämne  
Här kan du välja det datafält, vars innehåll ska infogas som ämne i dialogrutan Egenskaper.  
Filnamn för mallen  
I det här området definieras namn för och ev. beskrivning av dokumentmallen.  
Namn  
I det här textfältet kan du definiera dokumentmallens namn.  
Info  
Här kan du mata in texten som ska infogas som dokumentinfomation för den nya dokumentmallen i fältet Beskrivning i dialogrutan Egenskaper.  
Filnamn  
Här bestämmer du hur filnamnet för det skapade dokumentet ska börja.  
Automatiskt  
Markera den här rutan om %PRODUCTNAME ska använda filnamnet automatiskt.  
Prefix  
Texten under Prefix föreslås som filnamn för det skapade dokumentet.  
Du kan ändra texten i textfältet.  
Målkatalog...  
När du klickar på den här kommandoknappen öppnas dialogrutan Välj ut sökväg, där du kan ange var det skapade dokumentet ska arkiveras.  
Gå vidare till AutoPilot Brev - sida 9  
Gå vidare till AutoPilot Fax - sida 8  
Gå vidare till AutoPilot PM - sida 5  
Gå vidare till AutoPilot Agenda - sida 6  
AutoPilot Brev - sida 9  
I det sista steget bestämmer du slutligen om logotyp och avsändare ska upprepas på de följande sidorna i dokumentet och från vilka pappersfack (om skrivaren erbjuder detta alternativ) sidorna ska hämtas.  
Logotyp  
Här anger du på nytt på vilka sidor din logotyp ska visas.  
Alltid, Första sidan, Följande sidor, Skriv inte ut.  
Avsändare  
Här anger du på nytt på vilka sidor avsändaren ska visas.  
Alltid, Första sidan, Följande sidor, Skriv inte ut.  
Till sist anger du pappersmagasin.  
Om din skrivare stöder denna funktion, kan du här välja från vilka pappersmagasin den första sidan och de följande sidorna ska hämtas.  
Du kan t.ex. använda företagets papper till den första sidan och papper utan tryck till de följande sidorna.  
Första sidan  
Här bestämmer du från vilket pappersmagasin papperet till den första sidan i brevet ska hämtas.  
Följande sidor  
Här bestämmer du från vilket pappersmagasin papperet ska hämtas för sidan 2 och följande sidor.  
Ställ in...  
Om du trycker på den här kommandoknappen så visas dialogrutan Ställ in skrivare.  
AutoPilot Fax  
Med det här kommando öppnar du AutoPiloten för att skapa ett fax.  
Dessa kan du sedan skicka direkt via ett anslutet faxmodem (om sådant finns).  
%PRODUCTNAME har en mall för faxdokument som du kan anpassa efter din personliga smak med hjälp av AutoPiloten.  
AutoPiloten leder dig steg för steg genom de olika layoutelementen i dokumentmallen och ger dig möjlighet att välja mellan olika alternativ i varje steg.  
Den förminskade förhandsvisningen i dialogrutan ger dig ett intryck av vilken effekt de aktuella inställningarna har.  
I dialogrutan kan du när som helst ångra ett val eller hoppa över enskilda steg.  
Om du hoppar över ett steg använder AutoPiloten de aktuella förinställningarna.  
AutoPilot Fax - sida 2  
AutoPilot Fax - sida 6  
AutoPilot Fax - sida 7  
<<Tillbaka  
Med det här kommandot ser du alternativen som du valde i föregående steg.  
Kommandoknappen kan väljas från och med steg två.  
Nästa>>  
AutoPiloten använder de aktuella inställningarna i dialogrutan och går vidare till nästa steg.  
Om du har kommit till sista steget i dialogrutan går det inte att välja den här kommandoknappen.  
Färdigställ  
AutoPiloten skapar en ny dokumentmall enligt dina inställningar och sparar den på hårddisken.  
Med utgångspunkt från den nya dokumentmallen skapar %PRODUCTNAME ett nytt dokument med namnet "namnlösX" (X står för ett löpnummer) och visar det i arbetsområdet.  
%PRODUCTNAME sparar de aktuella inställningarna i AutoPiloten för den använda malltypen och använder dem som förinställningar nästa gång AutoPiloten öppnas.  
AutoPilot Fax - sida 1  
På den här sidan definierar du stil, rubrik och format för ditt faxdokument.  
Vilken stil vill Du använda?  
Välj en av följande stilar för faxet:  
Modern, Klassisk eller Elegant.  
Modern  
Här används främst sansserif-teckensnitt (utan seriffer).  
Klassisk  
Här används främst icke-proportionella teckensnitt.  
Elegant  
Här används främst antikvateckensnitt (med seriffer).  
Ange faxrubrik  
Här anger du texten som ska visas som överskrift i stor teckenstorlek uppe till vänster på faxet.  
Du kan även välja en överskrift bland några standardöverskrifter.  
Välj format för ditt fax  
Här kan du välja bland standardformaten som stöds av faxdrivrutinen.  
Gå vidare till AutoPilot Fax - sida 2  
AutoPilot Fax - sida 3  
På sida 3 i dialogrutan AutoPilot anger du avsändaren.  
Ange avsändaren  
Här anger du den avsändare som ska visas på samtliga fax som skapas med den här mallen.  
Avsändare  
I det här textfältet anger Du avsändare.  
Telefon  
Här kan du ange ditt telefonnummer.  
Telefax  
Här kan du ange ditt telefaxnummer.  
Uppdatera adress från användardata  
När du klickar på den här symbolen ersätts texten i avsändarfältet med en standardtext för avsändaren som hämtas från användardata.  
Position och storlek  
Här väljer du position och storlek för avsändarfältet på faxmallen.  
Välj position genom att klicka på dem.  
Du kan ställa in fältets storlek med rotationsfälten.  
Uppe till vänster  
Här placeras avsändarfältet uppe till vänster ovanför mottagaren.  
Uppe till höger  
Här placeras avsändarfältet uppe till höger bredvid mottagaren.  
Bredd  
Här kan du ställa in bredden för avsändarfältet.  
Höjd  
Här kan du ställa in höjden för avsändarfältet.  
Gå vidare till AutoPilot Fax - sida 4  
AutoPilot Fax - sida 4  
På den här dialogsidan anger du mottagaren.  
Databas  
Här väljer du den databas som innehåller poster med uppgifter för mottagaren.  
Databas  
Här väljer du tabellen från den markerade databasen där mottagaruppgifterna ska hämtas.  
Posterna i den här listrutan ändras beroende på vad du väljer i den vänstra listrutan Databas.  
Telefon  
Välj databasfältet, vars innehåll ska infogas som mottagarens telefonnummer i mallen.  
Telefax  
Välj databasfältet, vars innehåll ska infogas som mottagarens telefaxnummer i mallen.  
Adress  
Här kan du mata in mottagarens adress och / eller sammanställa den från databasfälten.  
Det senare alternativet är lämpligt för standardfax (kopplad utskrift).  
Databasfält  
Du kan infoga dem i adressfältet genom att klicka på dem med musen.  
Pil till vänster  
Det infogas där markören står i adressfältet.  
Styckebrytning  
Klicka här om du vill infoga en styckebrytning där markören står i adressfältet.  
Gå vidare till AutoPilot Fax - sida 5  
AutoPilot Fax - sida 5  
På sidan 5 bestämmer du vilka element faxet ska innehålla, t.ex. datum, ärenderad o.s.v.  
Vilka element skall Ditt fax innehålla?  
Här bestämmer du om olika element som brukar finnas i affärsfax ska användas i din mall.  
Datum  
Markera den här rutan om du vill infoga aktuellt datum (hämtas från operativsystemet) i faxet.  
Datum  
Här väljer du datumformat.  
Klockslag  
Markera den här rutan om du vill infoga aktuellt klockslag (hämtas från operativsystemet) i faxet.  
Klockslag  
Här väljer du klockslagets format.  
Ärenderad  
Markera den här rutan om du vill infoga en ärenderad i faxet.  
Ärenderad  
Här skriver du ärenderadens text.  
Kopia till  
Markera den här rutan om texten Kopia till ska infogas i faxet.  
1.  
För information  
Markera den här rutan om du vill infoga standardtexten För information i faxet.  
För information  
Använd standardtexten eller redigera den enligt dina önskemål.  
2.  
Att göra  
Om du markerar den här rutan infogas standardtexten Att göra i faxet.  
Att göra  
Använd standardtexten Att göra eller ändra den.  
3.  
Kommentera  
Markera den här rutan om du vill infoga denna standardtext i faxet.  
Kommentera  
Använd standardtexten i faxet eller redigera den enligt dina önskemål.  
4.  
Tack för lånet!  
Markera den här rutan om du vill infoga denna standardtext i faxet.  
Tack för lånet!  
Infoga texten i faxet eller redigera den.  
Fortsätt till AutoPilot Fax - sida 6  
AutoPilot Fax - sida 8  
På sidan 8 talar AutoPiloten om att du har gjort alla inställningar som behövs för den nya faxmallen.  
Klicka på Färdigställ så skapar %PRODUCTNAME faxmallen åt dig.  
AutoPilot PM  
Med det här kommandot startar du AutoPiloten för att skapa ett PM.  
Den hjälper dig att utforma dokumentmallar för PM.  
%PRODUCTNAME levereras med en mall för PM, som Du med hjälp av AutoPiloten kan anpassa till Dina personliga behov.  
AutoPiloten vägleder Dig steg för steg genom de olika elementen i dokumentmallen, och för varje redigeringssteg har Du olika alternativ att välja mellan.  
I dialogrutan finns en liten ruta för förhandsvisning som ger Dig en uppfattning om hur inställningarna påverkar resultatet.  
Du kan när som helst under processen ångra ett visst val; och Du kan också hoppa över enskilda redigeringssteg.  
Om Du hoppar över ett steg, använder AutoPiloten det stegets aktuella inställningar.  
AutoPilot PM - sidan 4  
<<Tillbaka  
De inställningar som Du just har gjort behålls.  
Den här kommandoknappen kan förstås inte användas vid det första redigeringssteget.  
Nästa>>  
AutoPiloten sparar inställningarna i den dialogruta som är öppen och går till nästa redigeringssteg.  
Om Du har kommit till den sista dialogrutan kan knappen förstås inte användas.  
Färdigställ  
AutoPiloten skapar på basis av de val Du har gjort en ny dokumentmall och sparar den på hårddisken.  
Med utgångspunkt från den nya dokumentmallen skapar %PRODUCTNAME ett nytt dokument med namnet "namnlös X" (X står för ett löpnummer) och visar detta i arbetsområdet.  
De aktuella inställningarna för den använda malltypen i AutoPiloten sparas och används som mall nästa gång Du använder AutoPiloten.  
AutoPilot PM - sida 1  
På dialogrutans första sidan definierar du vilken stil ditt PM ska skapas med.  
Dessutom bestämmer du vilken rubrik PM:et ska ha och om rubriken ska ersättas av ett grafikobjekt.  
Vilken stil vill Du använda?  
Välj en stil för ditt PM här:  
Modern, Klassisk eller Elegant.  
Modern  
Här används främst sanserif-teckensnitt (utan seriffer).  
Klassiskt  
Här används främst icke-proportionella teckensnitt.  
Elegant  
Här används främst antikvateckensnitt (med seriffer).  
Ange rubrik för Ditt PM  
Här anger du om PM:ets rubrik ska bestå av en text eller ett grafikobjekt.  
Som text  
Klicka här för att definiera en text som PM-rubrik.  
Som text  
Välj text bland standardtexterna i listrutan eller mata in en egen text.  
Som grafik  
Klicka på knappen Grafikurval när Du ska välja en grafikfil.  
Grafikurval...  
Med den här kommandoknappen öppnar du en dialogruta som liknar dialogrutan Infoga grafik.  
Gå vidare till AutoPilot PM - sida 2  
AutoPilot PM - sida 2  
Här bestämmer du vilka standardelement som ska ingå i ditt PM: datum, ärenderad o.s.v.  
Vilka element skall Ditt PM innehålla?  
Här anger du vilka vanliga PM-element som ska ingå i PM-mallen.  
I förhandsvisningsfältet ser du hur elementen påverkar PM:ets utseende när de markeras.  
Datum  
Markera den här rutan om du vill infoga aktuellt datum (hämtas från operativsystemet) i ditt PM.  
Datum  
Här väljer du datumformat.  
Ärenderad  
Markera den här rutan om du vill visa en ärenderad.  
Ärenderad  
Skriv ärenderadens text här.  
Till  
Markera den här rutan om du vill infoga texten Till i PM:ets huvud.  
Kopia till  
Markera den här rutan om du vill infoga texten Kopia till i PM:ets huvud.  
Från  
Markera den här rutan om du vill infoga texten Från i PM:ets huvud.  
1.  
Prioritet  
Markera den här rutan om du vill infoga texten Prioritet i PM:ets huvud.  
Prioritet  
Använd standardtexten eller redigera den enligt dina önskemål.  
2.  
Att göra tills  
Om ditt PM ska innehålla texten Att göra tills ska du markera den här rutan.  
Att göra tills  
Använd standardtexten eller redigera den enligt dina önskemål.  
3.  
Bilaga / or  
Markera den här rutan om texten Bilaga / or ska finnas i ditt PM.  
Bilaga / or  
Använd standardtexten eller redigera den enligt dina önskemål.  
4.  
Tom ruta  
Markera den här rutan om du vill infoga ytterligare text i PM:ets huvud.  
Tomt textfält  
Ange en text för ditt PM-element här.  
Gå vidare till AutoPilot PM - sida 3  
AutoPilot PM - sida 3  
På sidan 3 definierar du vilka element som ska visas på de följande sidorna i ett flersidigt PM.  
Vilka element vill Du placera i sidhuvudet på de följande sidorna?  
Här bestämmer du vilka vanliga PM-element som ska stå i sidhuvudet på de följande sidorna i PM:et.  
Datum  
Markera den här rutan om du vill att datum ska visas även på de följande sidorna.  
Den här rutan går bara att aktivera om du har valt datumvisning för första sidan i PM:et.  
Rubrik  
Markera den här rutan om du även vill infoga rubriken i sidhuvudet på de följande sidorna i ditt PM.  
Sidnummer  
Markera här för att sidnummer ska visas även på de följande sidorna.  
Skiljelinje mot text  
Markera den här rutan om du vill infoga en avgränsande linje mellan PM:ets huvud och texten.  
Vilka element vill Du placera i sidfoten på alla sidor?  
Här bestämmer du vilka vanliga PM-element som ska stå i sidfoten på samtliga sidor i PM:et.  
Datum  
Markera den här rutan om du vill att datum ska visas i sidfötterna.  
Den här rutan går bara att aktivera om du har valt datumvisning för första sidan i PM:et.  
Sekretessnivå  
Markera här för att infoga en anmärkning om sekretessnivån i sidfötterna.  
Sekretessnivå  
Skriv text här för en anmärkning om sekretessnivån.  
Nästa sidnummer  
Markera här om du vill att sidfoten ska innehålla information om antal efterföljande sidor.  
Skiljelinje för text  
Markera den här rutan om du vill infoga en avgränsande linje mellan text och sidfot.  
Gå vidare till AutoPilot PM - sida 4  
AutoPilot PM - sida 5  
På sidan 8 talar AutoPiloten om att du har gjort alla inställningar som behövs för den nya PM-mallen.  
Klicka på Färdigställ så skapar %PRODUCTNAME mallen åt dig och öppnar ett dokument som baserar på den nya mallen.  
AutoPilot Agenda  
Med det här kommandot får Du upp AutoPiloten för att skapa dagordningar.  
Den hjälper Dig att skapa dokumentmallar för dagordningar.  
Med den typen av dokument kan Du t ex skapa listor av dagordningstyp som kan användas för tal, möten o d.  
%PRODUCTNAME levereras med en mall för dagordningar, som Du med hjälp av AutoPiloten kan anpassa till Dina personliga behov.  
AutoPiloten vägleder Dig steg för steg genom de olika elementen i dokumentmallen, och för varje redigeringssteg har Du olika alternativ att välja mellan.  
Den förminskade förhandsvisningen i dialogrutan ger dig möjlighet att se effekten av de aktuella inställningarna.  
I dialogrutan kan du när som helst ångra ett val eller hoppa över enskilda steg.  
Om Du hoppar över ett steg, använder AutoPiloten det stegets aktuella inställningar.  
AutoPilot Agenda - sidan 5  
<<Tillbaka  
Dialogrutan återgår till valmöjligheterna i föregående redigeringssteg.  
De inställningar som Du just har gjort behålls.  
Kommandoknappen kan inte väljas förrän du har nått det andra steget.  
Nästa>>  
AutoPiloten använder de aktuella inställningarna i dialogrutan och övergår till nästa redigeringssteg.  
Om Du har kommit till den sista dialogrutan kan knappen förstås inte användas.  
Färdigställ  
AutoPiloten skapar en dokumentmall baserad på Dina inställningar och sparar denna på hårddisken.  
Med utgångspunkt från den nya dokumentmallen skapar %PRODUCTNAME ett nytt dokument med namnet "namnlös X" (X står för ett löpnummer) och visar detta i arbetsområdet.  
De aktuella inställningarna i AutoPiloten för den använda malltypen sparas och används som mall nästa gång Du använder AutoPiloten.  
AutoPilot Agenda - sida 1  
Här väljer du stil för dagordningen och anger rubrik.  
Alternativt kan du lägga in ett grafikobjekt i rubriken.  
Vilken stil vill Du använda?  
Här väljer du stil för mallen:  
Modern, Klassisk eller Elegant.  
Modern  
Här används främst sanserif-teckensnitt (utan seriffer).  
Klassisk  
Här används främst icke-proportionella teckensnitt.  
Elegant  
Här används främst antikvateckensnitt (med seriffer).  
Ange rubrik för mötet  
Här anger du den rubrik som ska visas på dagordningen.  
Logotyp  
Markera den här rutan om du vill använda en logotyp.  
Klicka på Grafikurval och välj en grafikfil i den dialogruta som visas.  
Grafikurval...  
Med den här kommandoknappen öppnar du dialogrutan Välj logotyp.  
Gå vidare till AutoPilot Agenda - sida 2  
AutoPilot Agenda - sida 2  
Här anger du datum, tidpunkt och plats för mötet.  
Ange datum och tid för mötet  
Ange datum och tidpunkt i dessa rotationsfält.  
Datum  
Ange datum för mötet här.  
Tidpunkt  
Här anger du klockslaget då mötet börjar.  
Ange plats för mötet  
I det här textfältet anger du var mötet äger rum.  
Vilka alternativ skall agendan innehålla?  
Här markerar du de rutor vars text ska infogas som alternativ i dagordningens huvud.  
Anledning  
Markera den här rutan om texten Anledning ska finnas i huvudet på dagordningen.  
Ta med  
Markera den här rutan om texten Ta med ska finnas i huvudet på dagordningen.  
Förbered  
Markera den här rutan om texten Förbered ska finnas i huvudet på dagordningen.  
Anmärkningar  
Markera den här rutan om texten Anmärkningar ska finnas i huvudet på dagordningen.  
Gå vidare till AutoPilot Agenda - sida 3  
AutoPilot Agenda - sida 3  
På sidan 3 väljer du vilka namn som ska finnas på med dagordningen.  
Vilka namn skall agendan innehålla?  
Här markerar du rutorna för namnen som ska finnas med i dagordningens huvud.  
Du kan välja bland "Kallat av", "Ledning", "Protokoll", "Deltagare", "Inbjudna", "Experter" och "Utvärdering ".  
Gå vidare till AutoPilot Agenda - sida 4  
AutoPilot Agenda - sida 4  
På den här sidan i dialogrutan anger du punkterna på dagordningen.  
Dialogrutan innehåller flera rader för dagordningspunkter.  
Först visas sex rader, men du kan öppna fler rader med hjälp av pilknappen.  
Mata in text för varje punkt som du vill ha med på dagordningen i textfältet Dagordningspunkt.  
Du kan dessutom ange en ansvarig.  
Ange tid i minuter för dagordningspunkten i rotationsfältet Tidslängd.  
Dagordningspunkt  
Här skriver du en text för dagordningspunktens rubrik.  
Ansvarig  
Här anger du namnet på den ansvarige.  
Tidslängd  
Här anger du planerad tidsåtgång i minuter för dagordningspunkten.  
Gå vidare till AutoPilot Agenda - sida 5  
AutoPilot Agenda - sida 6  
I det sista steget väljer du om du behöver ett protokollformulär.  
Sedan visas meddelandet att all information som krävs för att skapa agendamallen har sammanställts.  
Klicka på Färdigställ för att skapa mallen och automatiskt öppna ett dokument som baseras på mallen.  
Vill Du använda ett protokollformulär för att dokumentera Ditt möte?  
Här kan du avslutningsvis välja om du vill använda ett protokollformulär.  
I formuläret kan du under mötets gång anteckna punkter som ska åtgärdas, vem som är ansvarig och när punkten ska vara åtgärdad.  
AutoPilot Presentation  
Med hjälp av AutoPiloten skapar du en presentation interaktivt.  
De presentationsmallar som medföljer %PRODUCTNAME kan du anpassa till din personliga smak med hjälp av AutoPiloten.  
AutoPiloten leder dig steg för steg genom de olika layoutelementen och för varje redigeringssteg har du olika alternativ att välja bland.  
AutoPilot Presentation startas automatiskt när du öppnar en ny presentation via menyn Arkiv - Nytt.  
Du kan hindra AutoPiloten från att starta automatiskt genom att markera rutan Visa inte den här dialogrutan mer på första sidan.  
Du får samma effekt, om du, under Verktyg - Alternativ - Presentation - Allmänt, avmarkerar alternativet Starta med AutoPiloten.  
I varje dialogruta kan du när som helst ångra ett val eller hoppa över enskilda steg.  
Om du hoppar över ett steg, använder AutoPiloten de aktuella förinställningarna.  
<< Tillbaka  
Genom att klicka på den här kommandoknappen återgår du till föregående arbetssteg.  
De aktuella inställningarna bibehålls.  
Den här knappen går bara att använda fr.o.m. det andra redigeringssteget.  
Nästa >>  
AutoPiloten använder dina inställningar och går till nästa sida.  
När du har kommit till det sista steget i dialogrutan kan du inte välja den här kommandoknappen.  
Färdigställ  
Du kan sedan spara mallen med vilket namn du vill.  
%PRODUCTNAME Impress sparar de aktuella inställningarna i AutoPiloten och använder dessa som standard nästa gång AutoPiloten öppnas.  
AutoPilot Presentation - sida 1  
På den första sidan definierar du typ av presentation och väljer en tillhörande mall.  
Typ  
Här bestämmer du typ av presentation.  
Tom presentation  
Välj det här alternativfältet om du vill skapa en ny, tom presentation.  
Från mall  
Med det här alternativet öppnar du en listruta där du kan välja bland ett stort antal redigerbara presentationsmallar.  
Öppna en redan befintlig presentation  
Om du redan sparat några presentationer och väljer det här alternativet öppnas en lista över presentationerna.  
Om du vill ladda en presentation som finns på annat ställe på hårddisken, dubbelklickar du på posten Annan position.  
Dialogrutan Öppna visas.  
Listrutor med alternativ (bara om du markerat "Från mall")  
I den övre rutan kan du välja om du vill ha förslag till presentationer, utbildning eller presentationsbakgrunder.  
I listrutan nedanför kan du välja en av mallarna genom att klicka på den.  
Listruta med alternativ (bara om du markerat "Öppna en redan befintlig presentation")  
Du kan välja en av presentationerna som visas här och fortsätta att redigera den i AutoPiloten.  
Via posten Annan position kommer du till dialogrutan Öppna där du kan öppna en presentation som sparats i en valfri katalog.  
Förhandsvisning  
I förhandsvisningsfönstret visas den mall du valt.  
Du aktiverar / stänger av förhandsvisningen genom att klicka i kryssrutan.  
Visa inte den här dialogen mer  
Om du aktiverar den här rutan startas AutoPiloten i fortsättningen bara om du uttryckligen väljer det via menyn Arkiv - AutoPilot - Presentation.  
På menyn Verktyg - Alternativ - Presentation - Allmänt, finns området Nytt dokument, där kryssrutan Starta med AutoPiloten har samma funktion.  
Den här rutan visas bara om du har valt att skapa en presentation via menyn Arkiv - Nytt - Presentation.  
Fortsättning följer på AutoPilot Presentation - sida 2.  
AutoPilot Presentation - sida 2  
På den andra sidan väljer du presentationsmedium och bakgrund för presentationen.  
Välj en sidformatmall  
Här kan du tilldela den presentation som du valde på sidan 1 i AutoPiloten en annan sidformatmall.  
I den övre rutan kan du välja bland tre sidformatmalltyper.  
I listrutan nedanför kan du välja en av mallarna och lägga till den till presentationen genom att klicka på den.  
Välj ett presentationsmedium  
Original  
Du väljer det här alternativet om du vill använda original-sidformatet från mallen.  
Overhead  
Välj det här alternativet om du vill skriva ut presentationen på overheadfilm.  
Papper  
Välj det här alternativet om du vill skriva ut presentationen på papper.  
Bildskärm  
Det här alternativet innebär en ren bildskärmspresentation.  
Alternativet Bildskärm är förinställt.  
Dia  
Om du vill använda diabilder som visningsmedium väljer du det här alternativet.  
Fortsättning följer på AutoPilot Presentation - sida 3.  
AutoPilot Presentation - sida 3  
På den här sidan bestämmer du vilken typ av presentation du ska göra.  
Välj en diabildsväxling  
I det här området kan du tilldela din presentation effekter och definiera deras hastighet.  
Effekt:  
Välj en lämplig effekt i listan och klicka på den för att använda den i presentationen.  
Hastighet:  
Här bestämmer du med vilken hastighet effekten ska fungera.  
Du kan välja mellan "Långsamt", "Medel" och "Fort ".  
Välj typ av presentation  
Här definierar du förloppet för hela presentationen.  
Om du ändrar dig senare kan du göra andra inställningar via menyn Presentation.  
Standard  
Om du väljer alternativet Standard utförs presentationen som helskärmsvisning med den hastighet du angett.  
Du växlar bild genom att klicka med musen eller trycka på en särskild tangent (t.ex. returtangenten).  
Automatisk  
Markera det här alternativfältet om du vill att bildskärmspresentationen ska löpa automatiskt och starta på nytt efter en definierad paus.  
I rotationsfälten kan du göra mera detaljerade inställningar.  
Tid per sida  
Här definierar du visningstiden för enskilda diabilder i presentationen.  
Paustid  
I det här fältet anger du hur lång paus det ska vara mellan de olika presentationssekvenserna.  
Visa logotyp  
Välj det här alternativet om du vill att %PRODUCTNAME -logotypen ska visas på paussidan mellan presentationssekvenserna.  
Fortsättning följer på AutoPilot Presentation - sida 4.  
Om du har valt "Tom presentation" på sida 1 avslutas AutoPiloten och du kan skapa en ny presentation med egna inställningar.  
AutoPilot Presentation - sida 4  
Här kan du ange ditt företags namn och temat för presentationen och dessutom formulera grundidéer för presentationen.  
Beskriv dina grundidéer  
Här kan du formulera och skriva in dina tankar.  
Vad är Ditt namn eller Ditt företags namn?  
Skriv in fitt namn eller företagets namn i det här textfältet.  
Vilket tema har Din presentation?  
Här anger du det tema som du har valt för presentationen.  
Fler idéer som borde nämnas?  
I det här fältet kan du skriva in ytterligare idéer eller mål som du vill ta med i presentationen.  
Fortsättning följer på AutoPilot Presentation - sida 5.  
AutoPilot Presentation - sidan 5  
Här kan du bestämma vilka sidor som AutoPiloten ska ta med i presentationen.  
Välj de önskade sidorna  
I listrutan i det här området visas alla sidor som hör till den presentationsmall som du har valt.  
Genom att klicka på en sida infogar du den eller tar bort den från dokumentet.  
Om du klickar på det lilla plustecknet framför sidornas namn visas tillhörande underordnade punkter.  
Dina val visas i förhandsvisningsfönstret om du har markerat Förhandsvisning.  
Skapa sammanfattning  
Markera den här rutan om du vill skapa en sammanfattning av allt presentationsinnehåll.  
Tillbaka till huvudsidan för Autopilot Presentation....  
AutoPilot för webbsida  
Med det här kommandot startar du AutoPiloten för att skapa en webbsida.  
Vilken mall ska användas?  
Välj en mall för din webbsida i den här listrutan.  
Beroende på vilken mall du väljer fylls webbsidan med olika objekt på olika positioner.  
Du kan flytta, redigera och radera objekten på webbsidan.  
Vilken stil ska användas?  
Välj en stil för din webbsida i den här listrutan.  
Allt efter stil byts färger, bakgrund, teckensnitt, punkter och linjer.  
Skapa mall  
Den här rutan behöver du om du vill spara webbsidan som dokumentmall när du har skapat den med AutoPilot.  
Markera rutan innan du klickar på Färdigställ.  
I dialogrutan Dokumentmallar definierar du ett namn samt den kategori där den nya mallen ska sparas.  
I fortsättningen har du tillgång till den via menyn Arkiv - Nytt - Mallar och dokument.  
Du kan omvandla vilket som helst av dina öppnade dokument till en mall i efterhand.  
Med menyn Arkiv - Dokumentmall - Spara öppnar du dialogrutan Dokumentmallar, där du anger de uppgifter som behövs.  
Färdigställ  
Klicka på denna kommandoknapp för att färdigställa webbsidan med de aktuella inställningarna.  
Avbryt  
Om du stänger dialogrutan med kommandoknappen Avbryt, raderas den nya webbsidan.  
När AutoPilot har avslutats och den skapade webbsidan sparas för första gången, kopieras de använda grafiska objekten till den katalog där även filen har sparats.  
Samma sak sker om ett dokument sparas för första gången och dokumentet har skapats av en mall som genererats med AutoPilot.  
De grafiska objekten som finns i mallarna i AutoPilot kommer från Gallery i %PRODUCTNAME.  
När du sparar, kopieras dessa till den nya katalogen och sökvägarna i filen anpassas på motsvarande sätt.  
Autopilot - Formulär  
Med det här kommandot startar du AutoPiloten för att skapa ett formulär.  
Du väljer egenskaperna för formuläret på följande sätt:  
AutoPilot formulär:  
Databasurval  
På den här sidan i AutoPiloten bestämmer du för vilken tabell eller sökning du vill skapa ett formulär och vilka fält som du vill använda i formuläret.  
Datakälla  
Välj ut datakällan som du vill skapa formuläret för.  
Tabeller eller sökningar  
Välj ut tabellen eller sökningen som ska ligga till grund för formuläret.  
Existerande fält  
I den här listrutan visas namnen på datafälten från databastabellen.  
Du kan markera ett fält i den vänstra listan genom att klicka på det, eller så kan du använda tangenterna Skift eller Kommando Ctrl om du vill markera flera fält.  
->  
Klicka här om du vill använda det eller de markerade datafälten för formuläret.  
=>>  
Klicka här om du vill använda alla visade datafält för formuläret.  
< -  
Klicka här om du vill ta bort det eller de markerade datafälten från den högra listan.  
Det visas sedan i den vänstra listan igen.  
<<=  
Om du klickar här tas alla datafält som du har valt ut för formuläret tillbaka igen.  
Fält i formulär  
Här ser du de datafält som används i formuläret.  
Visning av binära fält  
Här väljer du hur binära fält ska behandlas i formuläret.  
Binära fält som grafik  
Om du väljer det här alternativet används binära fält som grafik i formuläret.  
Ignorera binära fält  
Om du väljer det här alternativet används inte binära fält i fomuläret.  
Gå vidare till AutoPilot formulär - Utformning  
AutoPilot formulär:  
Utformning  
På den här sidan i AutoPiloten väljer du en stil för det skapade formuläret.  
Dokumentet visar de olika ändringarna direkt utan att du måste stänga AutoPiloten först.  
Placering av DB-fält  
I kolumner - etiketter till vänster  
Markera det här alternativet om datafälten ska placeras kolumnorienterat.  
I kolumner - etiketter uppe  
Markera det här alternativet om datafälten ska placeras optimerat.  
Som tabell  
Markera det här alternativet om datafälten ska placeras i tabellform.  
Marginaljusterat - etiketter till vänster  
Markera det här alternativet om du vill att rubrik och data ska placeras bredvid varandra.  
Marginaljusterat - etiketter uppe  
Markera det här alternativet om du vill att rubrik och data ska placeras ovanför varandra.  
Fältinramning  
Utan inramning  
Fälten får ingen kant.  
3D-look  
Fälten visas i en 3D-look.  
Flat  
Fälten visas flata.  
Sidformatmallar  
Välj en av mallarna i listrutan för det nya formuläret.  
Justering av etikettfält  
Vänsterjusterat  
Etiketterna vänsterjusteras.  
Högerjusterat  
Etiketterna högerjusteras.  
Bakgrundsbild  
Sida vid sida  
Bakgrundsbilden visas sida vid sida.  
Skalat  
Bakgrundsbilden visas skalat.  
HTML-export  
Den här AutoPiloten hjälper dig att publicera dina %PRODUCTNAME Draw - eller %PRODUCTNAME Impress-dokument i HTML-format.  
När du exporterar flersidiga dokument underlättar den här AutoPiloten arbetet avsevärt.  
Du får bl.a. en automatiskt skapad översiktssida och, om du vill, ramar, navigationselement och andra hjälpelement.  
Olika fortsättningssidor visas beroende på vilka val du gör på den andra sidan i AutoPiloten.  
<< Tillbaka  
Du kan gå tillbaka och se vilka val Du har gjort på föregående sida.  
Aktuella inställningar bibehålls.  
Denna knapp är endast tillgänglig fr o m det andra redigeringssteget.  
Nästa >>  
När Du klickar på den här knappen använder AutoPiloten de aktuella inställningarna i dialogrutan och går vidare till nästa sida.  
Om Du har kommit till den sista sidan i dialogrutan kan knappen inte väljas.  
Färdigställ  
AutoPiloten skapar nya dokument baserade på dina inställningar och sparar dem på hårddisken.  
%PRODUCTNAME sparar de aktuella inställningarna i AutoPiloten och använder dem som förinställningar nästa gång AutoPiloten öppnas.  
HTML-export - sida 1  
På den första sidan väljer du en färdig design eller skapar en ny design.  
De inställningar som du har valt för en export sparas automatiskt som design för andra exporter.  
Du kan ge designen ett namn i en liten dialogruta när du har klickat på Färdigställ.  
Tilldela design  
I det här området kan du börja skapa en ny design eller välja eller radera en befintlig.  
Någon exportfil raderas inte.  
Ny design  
Markera det här alternativet om Du vill definiera en ny design på Autopilotens följande sidor.  
Existerande design  
Markera det här alternativet om Du vill ladda en befintlig design från designlistan och använda den som utgångspunkt på de följande sidorna i Autopiloten.  
Designlista  
På den här listan ser Du de designer som Du redan har definierat.  
Radera markerad design  
Klicka på den här knappen när Du vill radera den design som Du har markerat på designlistan.  
HTML-export - sida 2  
På den här sidan väljer du typ av publicering.  
Du bestämmer bl.a. om ramar ska användas, om en titelsida ska skapas med och om de anteckningar som du har gjort till presentationssidor också ska visas.  
Typ av publicering  
I det här området gör du grundinställningar (t.ex. Skapa titelsida) för den kommande exporten.  
Standard-HTML-format  
Markera det här alternativet om de exporterade sidorna ska skapas som enkla HTML-sidor.  
Standard-HTML med ramar  
Markera det här alternativet om du vill skapa ramar.  
Den exporterade sidan skapas i huvudramen, medan en innehållsförteckning i form av hyperlänkar visas i en sidoram.  
Skapa titelsida  
Om du markerar den här kryssrutan skapas som inledning en titelsida.  
Visa anteckningar  
Om de anteckningar som hör till objektet också ska visas, markerar du den här rutan.  
Automatisk  
Tidsintervallen är de tider som du har definierat som visningstid för de olika diabilderna eller en och samma tid för alla diabilder.  
Som angivet i dokumentet  
Sidväxlingen görs efter det tidsintervall som Du har angett för varje diabild i presentationen.  
Om Du har angett manuell sidväxling, inväntar HTML-presentationen en tangenttryckning.  
Automatisk  
Sidväxlingen görs automatiskt efter en fastställd tid, oavsett vilka tider som har angetts i presentationen.  
Tid per sida  
Här väljer du den tid per sida som varje diabild ska visas.  
Kontinuerlig  
Om du markerar rutan Kontinuerlig, börjar HTML-presentationen om med den första bilden när den sista har visats.  
WebCast  
Vid WebCast-export genereras automatiskt skript för webb-servrar som stöder Perl eller ASP.  
En föredragshållare (t ex i en presskonferens över telefon med beledsagande bildvisning över Internet) kan på så sätt växla sidorna i åskådarens webbläsare.  
Mer information om WebCast-export finns längre ned.  
Active Server Page (ASP)  
Med det här alternativet skapar Du ASP-sidor för WebCast-exporten.  
Den HTML-presentation som Du skapar på detta sätt kan bara förmedlas av en webbserver som stöder ASP.  
Perl  
Med det här alternativet skapar Du HTML-sidor och Perl-skript för WebCast-exporten.  
URL för åhörare  
Här anger Du den URL-adress (absolut eller relativ) som den som ska titta på presentationen i sin webbläsare måste ange för att kunna se presentationen.  
URL för presentation  
Här anger Du den URL-adress (absolut eller relativ) under vilken den HTML-presentation som Du har skapat lagras på webbservern.  
URL för perl-skript  
Här anger Du URL-adressen för perl-skripten.  
Även denna URL kan vara absolut eller relativ.  
Närmare information om WebCast-export  
Active Server Pages (ASP) och Perl.  
För WebCast behövs åtminstone en HTTP-server som stöder antingen Perl eller ASP som scripting.  
Vilken variant av exporten Du väljer beror således främst på den HTTP-server som Du använder.  
Dessutom måste Du ha solida kunskaper om hur man använder webbservern och ASP respektive Perl, så att Du kan arbeta vidare med de filer som skapats av WebCast-exporten.  
WebCast via ASP  
Exporten  
För export enligt ASP väljer du i ett öppet %PRODUCTNAME Impress-dokument menykommandot Arkiv - Exportera Dialogrutan Exportera visas där du kan välja Webbsida som filtyp.  
När du har valt en katalog och angett ett filnamn klickar du på Spara.  
Vid export som ASP bör du ge HTML-filen ett "hemligt" filnamn, se vidare nedan.  
Nu visas dialogrutan HTML-export.  
Den skriver in ett antal filer i den valda katalogen.  
Det angivna filnamnet kommer senare att användas av föredragshållaren för att växla sidorna hos åhöraren.  
Som mapp kan Du välja en mapp eller en HTTP-URL-adress på HTTP-servern.  
Du kan också överföra de filer Du har skapat till HTTP-servern senare, t ex via FTP.  
Observera att WebCast bara fungerar om filerna hämtas från HTTP-servern.  
En allmän regel vid HTML-export är att Du måste exportera olika dokument i olika mappar.  
Det går inte att göra två HTML-exporter i samma mapp, eftersom den andra exporten delvis skulle skriva över den första.  
Välj WebCast som publiceringstyp på sidan 2 i autopiloten för HTML-export.  
I det alternativområde för WebCast som då visas markerar Du Active Server Pages (ASP).  
Nu kan Du göra ytterligare inställningar eller starta exporten med kommandoknappen Slutför.  
Användning  
Så snart de exporterade filerna är tillgängliga på en HTTP-server, kan Du använda WebCast-tekniken.  
Exempel  
Du har installerat Microsoft Internet Information Server på datorn.  
Som startträd för Dina HTML-dokument har Du vid installationen angett mappen C:\Inet\wwwroot\foredrag.  
Datorns URL-adress bör vara http: / /minserver.com.  
De filer som skapades av exportfunktionen har Du sparat i mappen c:\Inet\wwwroot\foredrag\.  
I denna mapp skapar exportfunktionen en HTML-fil som t ex kan få filnamnet hemlig.htm.  
Du har angett detta namn i dialogrutan Spara (se ovan).  
Föredragshållaren kan nu ladda HTML-exporten i en valfri HTTP-läsare med stöd för JavaScript genom att skriva in URL-adressen http: / /minserver.com / foredrag / hemlig.htm.  
Via en serie av formulärfält kan han ändra den visade sidan.  
Ett valfritt antal åhörare kan nu via webbadressen http: / /minserver.com / föredrag / webcast.asp titta på den sida som föredragshållaren har valt.  
Via denna URL kan den aktuella sidan inte bytas.  
Om föredragshållaren hemlighåller den URL som han använder (därför namnförslaget hemlig.htm), kan föredraget inte saboteras.  
Du bör se till att HTTP-servern inte tillåter visning av mappar.  
WebCast via Perl  
Export  
I ett öppnat %PRODUCTNAME Impress-dokument exporterar du med menykommandot Arkiv - Exportera.  
Nu visas dialogrutan Exportera där du väljer Webbsida som filtyp.  
När du har valt en katalog och matat in ett filnamn klickar du på Spara.  
Nu visas AutoPilot för HTML-export.  
Den här exportfunktionen kommer att skriva flera filer i den just valda katalogen.  
Det inmatade filnamnet används senare av föredragshållaren för att byta åhörarnas sidor.  
Som mapp ska Du välja en tom mapp.  
I AutoPilot HTML-export väljer Du på andra sidan WebCast som typ av publicering.  
Nu visas ett område med alternativ för WebCast, där aktiverar Du Perl.  
I inmatningsfältet URL för åhörare anger Du det filnamn som HTML-dokumentet för åhörarna har.  
I inmatningsfältet URL för presentation ska URL-adressen till mappen för presentationen anges.  
I inmatningsfältet URL för perl-skript anger Du URL-adressen för den önskade CGI-skript-mappen.  
Nu kan Du göra fler inställningar eller starta exporten via kommandoknappen Färdigställ.  
Användning  
De filer som har skapats genom exporten måste nu först implanteras på HTTP-servern, vilken måste ha Perl-stöd.  
Eftersom det finns ett stort antal olika typer av HTTP-servrar med Perl-stöd kan detta inte automatiseras.  
Här följer en allmän beskrivning av de arbetsmoment som behöver utföras.  
Se efter i handboken till servern eller fråga nätverksadministratören hur dessa arbetsmoment ska utföras på servern.  
Först måste de filer som har skapats vid exporten flyttas till de rätta mapparna på HTTP-servern.  
De filer som har filnamnstilläggen htm, jpg och gif läggs på HTTP-servern i den mapp vars URL-adress har angetts i inmatningsfältet URL för presentation.  
De filer som har filnamnstilläggen pl och txt läggs på HTTP-servern i den mapp vars URL-adress har angetts i inmatningsfältet URL för perl-skript.  
Denna mapp måste vara konfigurerad på ett sådant sätt att de perl-skript som ligger där verkligen utförs efter en HTTP-begäran.  
Under Unix-system är det nödvändigt att filer med filnamnstillägget pl även tilldelas motsvarande rättigheter som tillåter att de utförs av HTTP-servern.  
Detta görs i regel via kommandot chmod.  
Dessutom måste rättigheterna för filen currpic.txt vara så inställda att HTTP-servern kan skriva i denna fil.  
Nu bör Du kunna använda WebCast.  
Exempel  
Du har en Linux-dator med en installerad HTTP-server.  
Din HTTP-servers URL heter http: / /minserver.com.  
Utmapp för Dina HTML-dokument är mappen / /user / local / http /, Dina perl-skript finns i mappen / /user / local / http / cgi-bin /.  
Som filnamn vid exporten väljer Du hemlig.htm.  
Som URL för åhörare anger Du foredrag.htm.  
Som URL för presentation anger Du http: / /minserver.com / foredrag / och som URL för perl-skript väljer Du http: / /minserver.com / cgi-bin /.  
Ur den mapp som angetts vid exporten kopierar Du nu alla *.htm, *.jpg och *.gif-filer till mappen "/ /user / local / http / foredrag /" på Din HTTP-server.  
De filer som har filnamnstilläggen *.pl och *.txt kopierar Du till mappen "/ /user / local / http / cgi-bin /".  
Nu loggar Du in som root på servern och växlar till mappen '/ /user / local / http / cgi-bin /'.  
Med kommandot chmod kan Du ställa in de motsvarande rättigheterna.  
När Du är klar med installationen av perl-filerna, kan föredragshållaren leda föredraget under URL-adressen http: / /minserver.com / foredrag / hemlig.htm och åhörarna kan titta på föredraget under URL-adressen http: / /minserver.com / foredrag / foredrag.htm.  
HTML-export - sida 3  
På den här sidan väljer du grafiktyp och målbildskärmens upplösning.  
Spara grafik som  
I det här området definierar du formatet.  
Dessutom definierar du komprimeringsvärdet för exporten.  
GIF  
Markera här om du vill exportera sidorna som GIF-filer.  
GIF-filer är komprimerade, förlustfria och har maximalt 256 färger.  
JPG  
Markera här om du vill exportera sidorna som JPEG-filer.  
De kan innehålla fler än 256 färger.  
Komprimering  
Välj här komprimeringsfaktorn för JPEG-grafiken.  
Ett värde på 100% ger bästa kvalitet vid stora filer, medan en faktor på 25% ger de minsta filerna, men med sämre bildkvalitet.  
Bildskärmsupplösning  
Här bestämmer du upplösningen för målbildskärmen.  
Bilden matas ut med upp till 80% förminskning, beroende på vald upplösning.  
Låg upplösning (640x480 pixel)  
Välj låg upplösning när visningen ska vara relativt stor.  
Mediumupplösning (800x600 pixel)  
Välj mediumupplösning för en medelstor visning.  
Hög upplösning (1024x768 pixel)  
Välj en hög upplösning för en starkt förminskad visning.  
Exportera ljud vid sidväxling  
Om du markerar den här rutan, exporteras även ljudfiler som du har definierat som effekt vid sidväxling.  
HTML-export - sida 4  
På den här sidan anger du uppgifter som ska visas på den exporterade publikationens titelsida.  
Den här sidan hoppas över om du har avmarkerat kryssrutan Skapa titelsida eller om du har valt automatisk export eller WebCast-export.  
Information för titelsidan  
Om du på AutoPilotens andra sida har angett att du ska ha en titelsida, gör du motsvarande inmatningar här.  
Skapad av  
Ange här namnet på den som ska stå som publikationens författare.  
E-postadress  
Här anger du den e-postadress till vilken publikationens läsare kan skicka kommentarer eller frågor.  
Din hemsida  
Den infogas som hyperlänk i publikationen.  
Mer information  
I det här textfältet kan du föra in mer text som ska visas på titelsidan.  
Länk till kopia av originalpresentationen  
Om du vill infoga en länk till en kopia av originalet markerar du den här kryssrutan.  
HTML-export - sida 5  
På den här sidan i AutoPiloten väljer du en stil för kommandoknapparna för att navigera mellan publikationens sidor.  
Den här sidan hoppas över om du har avmarkerat kryssrutan Skapa titelsida eller om du har valt automatisk export eller WebCast-export.  
Välj ut stil för kommandoknappar  
Här anger Du om Du vill ha kommandoknappar i dokumentet och vilken stil de i så fall ska ha.  
Bara text  
Om du markerar den här rutan, infogas hyperlänkar bara som texter i stället för grafiska kommandoknappar.  
Urvalsfält  
Här kan Du välja mellan olika typer av grafiska kommandoknappar.  
HTML-export - sida 6  
På den sista sidan i AutoPiloten för HTML-export bestämmer du vilka färger publikationen ska ha.  
Formateringen av texterna hämtas från teckningen respektive presentationen.  
Sidan hoppas över om du har avmarkerat kryssrutan Skapa titelsida eller om du har valt automatisk export eller WebCast-export.  
Välj ut färgschema  
Här anger Du det färgschema och de färger som ska användas till text, bakgrund osv.  
Överta färgschema från dokument  
Om det här alternativet är markerat, övertas färgerna från den aktuella dokumentmallen.  
Använd browserfärger  
Om det här alternativet är markerat, används färginställningarna i läsarens webbläsare (browser).  
Använd eget färgschema:  
Med det här alternativet kan Du definiera egna färger för olika element i publikationen.  
Text  
Om Du klickar här kan Du välja färg på texten i publikationen i dialogrutan Färg.  
Hyperlänk  
Om Du klickar här kan Du välja färg på hyperlänkar i publikationen i dialogrutan Färg.  
Aktiv länk  
Om Du klickar här kan Du välja färg på aktiva hyperlänkar i publikationen i dialogrutan Färg.  
Använd länk  
Om Du klickar här kan Du välja färg på besökta hyperlänkar i publikationen i dialogrutan Färg.  
Bakgrund  
Om Du klickar på den här kommandoknappen öppnas dialogrutan Färg, där Du kan välja färg på publikationens bakgrund.  
AutoPilot för gruppelement  
AutoPilot för gruppelement startar automatiskt när du infogar en grupperingsram i ett dokument.  
Färdigställ  
Om du klickar här skapas objektet.  
Data  
På första sidan definierar Du vilka alternativfält gruppelementet ska innehålla.  
Vilka beteckningar skall alternativfälten få?  
Här anger Du separat för varje alternativfält dess beteckning.  
Överta  
>>  
Med denna kommandoknapp bekräftar Du alternativfältets namn och övertar det i listan Alternativfält.  
För varje alternativfält i gruppen som ska skapas anger du den önskade beteckningen och övertar det inmatade namnet till listan Alternativfält genom att klicka på pilknappen.  
Upprepa denna procedur tills alla alternativfält är definierade.  
Alternativfält  
Här listas alla alternativfält som ska tas med i gruppelementet.  
Ångra  
<<  
Med denna kommandoknapp kan Du ta bort ett redan definierat alternativfält.  
Markera den önskade posten innan Du klickar på kommandoknappen.  
AutoPilot för gruppelement:  
Standardfälturval  
Här anger du om ett visst alternativfält är förvalt.  
Den här standardinställningen antas om formuläret öppnas i användarläge. (Med den inställning som du gör här bestämmer du kontrollfältsegenskapen Standardstatus.)  
Skall ett alternativfält vara utvalt som standard?  
Här bestämmer Du om det ska finnas någon standardinställning för alternativgruppen.  
Ja, följande:  
Välj detta alternativ om något alternativfält ska vara aktivt som standard när formuläret öppnats.  
Det aktiva alternativfältet väljer Du i listrutan.  
Listruta  
Här väljer Du det alternativfält som ska vara aktivt som standard när formuläret öppnas.  
Här listas alla alternativfält som Du har definierat på den föregående sidan.  
Nej, inget fält skall vara utvalt  
Med detta alternativ kommer inget alternativfält att vara aktivt som standard.  
AutoPilot för gruppelement:  
Fältvärden  
Här kan du tilldela varje alternativfält ett referensvärde.  
Välj först ett fält i listan med alternativfält och skriv sedan in referensvärdet för detta fält.  
Vilket värde vill du tilldela varje alternativ?  
Här anger du ett tal eller en text som referensvärde.  
Alternativfält  
Markera här det alternativfält som ska tilldelas referensvärdet.  
AutoPilot för gruppelement:  
Databasfält  
Den här sidan visas om dokumentet är kopplat till en databas.  
Här anger du om referensvärdena ska sparas i databasen.  
Därför anger du här i vilket datafält referensvärdena ska sparas.  
Ett referensvärde kan i en databas representera gruppelementets aktuella status.  
Denna sida visas bara om dokumentet redan är kopplat till en databas.  
Vill du spara värdet i ett databasfält?  
Ja, i följande databasfält  
När Du väljer detta alternativ sparas referensvärdena i databasen.  
De skrivs i det datafält som Du väljer i listrutan.  
I listrutan finns alla fält i databasen som formuläret är kopplat till.  
Listruta  
Här väljer Du det datafält i vilket referensvärdena ska sparas.  
Nej, jag vill bara spara värdet i formuläret  
Med detta alternativ sparas referensvärdena inte i databasen utan bara i formuläret.  
AutoPilot för gruppelement:  
Skapa alternativgrupp  
På sista sidan anger du slutligen ett namn för alternativgruppen.  
Vilken beteckning skall din alternativgrupp ha?  
Ange den önskade beteckningen för alternativgruppen i textfältet.  
AutoPilot Dokumentkonverterare  
AutoPiloten konverterar dokument till XML-formatet som används av %PRODUCTNAME från och med version 6.0.  
AutoPiloten konverterar dokument och mallar från det binära formatet som %PRODUCTNAME använde innan version 6.0 samt dokument från Microsoft Word, Excel eller Powerpoint.  
Källfilerna läses bara och ändras alltså inte.  
Nya målfiler skrivs (med nytt filnamnstillägg), i samma eller en annan mapp.  
Dokumentkonverteraren omfattar följande sidor:  
Dokumentkonverterare Sammanfattning  
På den här sidan finns en sammanfattande text som informerar dig om vad som konverteras om du klickar på Konvertera.  
Dokumentkonverterare - första sidan  
På den här sidan definierar du om det är dokument från %PRODUCTNAME eller från Microsoft Office som ska konverteras och vilken dokumenttyp som ska konverteras.  
%PRODUCTNAME  
Välj det här alternativet om du vill konvertera binära %PRODUCTNAME -dokument (d.v.s. dokument som har skapats innan 6.0-versionen) till XML-dokument.  
Textdokument  
Markera den här rutan om du vill konvertera dokument i det gamla %PRODUCTNAME Writer-formatet *.sdw till *.sxw.  
Tabelldokument  
Markera den här rutan om du vill konvertera dokument i det gamla %PRODUCTNAME Calc-formatet *.sdc till *.sxc.  
Tecknings - / presentationsdokument  
Markera den här rutan om du vill konvertera dokument i det gamla %PRODUCTNAME Draw-formatet *.sda till *.sxd och %PRODUCTNAME Impress-formatet *.sdd till *.sxi.  
Samlingsdokument / formler  
Markera den här rutan om du vill konvertera dokument i det gamla %PRODUCTNAME Writer samlingsdokument-formatet *.sgl till *.sxg och %PRODUCTNAME Math-formatet *.smf till *.mml.  
Microsoft Office  
Välj det här alternativet om du vill konvertera Microsoft Office-dokument till %PRODUCTNAME -dokumentformatet XML.  
Word-dokument  
Markera den här rutan om du vill konvertera dokument i Microsoft Word-formatet *.doc till *.sxw.  
Excel-dokument  
Markera den här rutan om du vill konvertera dokument i Microsoft Excel-formatet *.xls till *.sxc.  
PowerPoint-dokument  
Markera den här rutan om du vill konvertera dokument i Microsoft PowerPoint-formatet *.ppt till *.sxi.  
Skapa loggfil  
Loggfilen visar vilka dokument som har konverterats.  
Här fortsätter du till nästa sida i dokumentkonverteraren  
Dokumentkonverterare - följande sidor  
På de här sidorna väljer du för varje malltyp och dokumenttyp från vilken mapp dokumentkonverteraren ska läsa och till vilken mapp den ska skriva.  
Mallar  
Här definierar du om och hur dokumentmallarna ska konverteras.  
Textmallar  
("Textmallar "står för den dokumenttyp som valdes på den föregående sidan i dokumentkonverteraren.)  
Markera den här rutan om du vill konvertera dokumentmallarna.  
inkl. underordnade kataloger  
Markera den här rutan om även de underordnade katalogerna till den valda mappen ska sökas igenom efter filer.  
Importera från  
Välj mappen som innehåller källfilerna.  
Spara i  
Välj mappen där målfilerna ska skrivas.  
...  
Den här kommandoknappen öppnar dialogrutan Välj ut sökväg.  
Dokument  
Här definierar du om och hur dokument ska konverteras.  
Textdokument  
("Textdokument "står för den dokumenttyp som valdes på den föregående sidan i dokumentkonverteraren.)  
Markera den här rutan om du vill konvertera dokumenten.  
Här kommer du tillbaka till AutoPilotens huvudsida Dokumentkonverterare  
AutoPilot Eurokonverterare  
Den här AutoPiloten hjälper dig att konvertera valutabelopp i %PRODUCTNAME Calc - och %PRODUCTNAME Writer-dokument till Euro.  
Om du konverterar filer får de inte vara öppna.  
Men det är också möjligt att använda eurokonverteraren på ett öppet %PRODUCTNAME Calc-dokument.  
I så fall visas dialogrutan som beskrivs i slutet av det här avsnittet.  
Observera att endast valuta från länder som infört euro som gemensam valuta konverteras.  
Omfattning  
Enskilt %PRODUCTNAME -dokument.  
Välj det här alternativet om bara en enda %PRODUCTNAME Calc - eller %PRODUCTNAME Writer-fil ska konverteras.  
Hela katalogen  
Välj det här alternativet om du vill att alla %PRODUCTNAME Calc - och %PRODUCTNAME Writer-dokument och mallar i en katalog ska konverteras.  
Valutor:  
Välj valutan som ska konverteras till euro här.  
Källkatalog / källdokument  
I det här textfältet anger du katalogen resp. namnet på filen (filerna) som ska konverteras.  
...  
Den här kommandoknappen öppnar en dialogruta där du kan hitta katalogen eller filen.  
Inklusive undermappar  
Aktivera den här rutan om du vill ta med alla underordnade mappar.  
Konvertera även fältkommandon och tabeller i textdokument  
Markera den här rutan om du förutom %PRODUCTNAME Calc-dokument även vill konvertera %PRODUCTNAME Writer-dokument.  
Upphäv tabellskydd temporärt utan säkerhetsfråga  
Om den här rutan är markerad upphävs tabellskyddet medan konverteringen pågår och återupprättas igen efteråt.  
Om tabellskyddet är försett med ett lösenord visas en dialogruta där du kan ange lösenordet.  
Målmapp  
Här anger du katalogen med sökväg där de konverterade filerna ska sparas.  
Här är redan den arbetskatalog förvald som har ställts in under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar - Arbetskatalog.  
...  
Med den här kommandoknappen öppnar du en dialogruta med vars hjälp du kan välja en katalog där de konverterade filerna ska placeras.  
Avbryt  
Klicka på den här kommandoknappen om Du vill stänga Eurokonverteraren.  
Hjälp  
Med den här kommandoknappen aktiverar du hjälpen till dialogrutan.  
Konvertera  
Här startar du konverteringen.  
Under konverteringen visas en sida med statusmeddelanden om hur konverteringen fortskrider.  
Tillbaka  
Från statussidan kommer du tillbaka till den första sidan i Eurokonverteraren med kommandoknappen Tillbaka.  
Om det aktuella dokumentet är ett %PRODUCTNAME Calc-dokument eller en mall, kan du starta Eurokonverteraren via en ikon på verktygslisten.  
Den här ikonen döljs enligt standardinställning; du ser den först när du visar den via kommandot Synliga knappar på verktygslistens snabbmeny.  
Eurokonverterare  
Dialogrutan Eurokonverterare visas med följande funktioner:  
Komplett dokument  
Markera det här fältet om Du vill att hela dokumentet ska konverteras.  
Valutor  
Välj valutan som ska konverteras till Euro i det här kombinationsfältet.  
Markering  
I det här området väljer du ut cellerna som ska konverteras om du inte har markerat Komplett dokument.  
Valutaområden till höger.  
I dokumentet visas det valda området som markering.  
När du vill konvertera klickar du på Konvertera.  
Cellmallar  
Alla celler med de valda cellmallarna konverteras.  
Valutaceller i det aktuella tabellarket  
Alla valutaceller i det aktuella tabellarket konverteras.  
Valutaceller i hela dokumentet  
Alla valutaceller i det aktuella dokumentet konverteras.  
Utvalt område  
Alla valutaceller konverteras som finns i ett område som har markerats innan konverteraren startades.  
Alla celler måste ha samma formatering för att de ska godtas som "Utvalt område".  
Mallar / Valutaområden  
Markera områdena som ska konverteras i listan.  
I dokumentet markeras de valda områdena så att du kan kontrollera dem.  
%PRODUCTNAME 5.2 databasimport  
Med det här kommandot startar du en AutoPilot som kan importera %PRODUCTNAME 5.2-databaser till %PRODUCTNAME %PRODUCTVERSION.  
Den här AutoPiloten ändrar, flyttar eller raderar inte dina länkar till databaser eller databasfiler som du har skapat i %PRODUCTNAME 5.2, t.ex. address.dbf.  
AutoPiloten använder informationen i *.sdb-filen i %PRODUCTNAME 5.2 och registrerar en ny datakälla i %PRODUCTNAME %PRODUCTVERSION.  
Uppgifterna är sedan tillgängliga i %PRODUCTNAME %PRODUCTVERSION, t.ex. under Verktyg - Datakällor eller i datakällvyn (F4).  
Den här AutoPiloten skapar inga kopior av tabeller.  
Det skapas t.ex. ingen kopia av en dbf-fil i dBase-format som ligger i din %PRODUCTNAME 5.2-katalog.  
Radera alltså inte dbf-filen!  
Om det finns sökningar eller formulär i den valda *.sdb-filen kan du ange i AutoPiloten att de ska läsas ut från *.sdb-filen och skapas som nya dokument i en katalog som du väljer.  
Färdigställ  
Det här kommandot skapar anslutningen av datakällan och stänger dialogrutan.  
%PRODUCTNAME 5.2 databasimport - Definiera källa  
Här väljer du databasfilen från %PRODUCTNAME 5.2 med tillägget *.sdb vars data du vill importera till %PRODUCTNAME %PRODUCTVERSION.  
Källa  
Ange sökvägen till en databasfil (*.sdb) från %PRODUCTNAME 5.2.  
Genomsök  
Här öppnar du en dialogruta där du kan leta efter en *.sdb-fil.  
Till nästa sida  
%PRODUCTNAME 5.2 databasimport - Element som ska importeras  
Här väljer du ut elementen som ska importeras.  
Mål  
Importera datakälla  
Markera den här rutan om du vill importera tabeller.  
Importera sökningar  
Markera den här rutan om du vill importera sökningar.  
Om du markerar rutan visas dialogrutan Formulärimport senare.  
Importera formulärdokument  
Markera den här rutan om du vill importera formulärdokument.  
Om du markerar rutan visas dialogrutan Sökningsimport senare.  
Till sidan Anpassa sÃ¶kvÃ¤g  
Till sidan FormulÃ¤rimport  
Till sidan SÃ¶kningsimport  
Till sidan Sammanfattning  
%PRODUCTNAME 5.2 databasimport - Anpassa sökväg  
Här anpassar du sökvägen till databasen.  
Den här sidan i AutoPiloten visas bara om du importerar en databas i *.dbf - eller textformat och det samtidigt finns en variabel i sökvägen till källdatabasen.  
Skriv den fullständiga sökvägen till källdatabasen utan att använda variablerna.  
Ny sökväg  
Ersätt variabeln i sökvägen med den fullständiga sökvägen.  
Till sidan Formulärimport  
Till sidan Sökningsimport  
Till sidan Sammanfattning  
%PRODUCTNAME 5.2 databasimport - Formulärimport  
Här väljer du ut formulären som ska importeras och deras målkatalog.  
Formulär  
Ange katalogen dit du vill kopiera formulären som dokument.  
Genomsök  
Här öppnar du en dialogruta där du kan välja katalog.  
formulär som ska importeras  
Här väljer du formulären som du vill kopiera som dokument.  
Alla  
Klicka här om du vill välja ut alla formulär.  
Inga  
Klicka här om du inte vill välja ut något formulär.  
Till sidan SÃ¶kningsimport  
Till sidan Sammanfattning  
%PRODUCTNAME 5.2 databasimport - Sökningsimport  
Här väljer du sökningarna som ska importeras och deras datakälla.  
Datakälla  
Ange datakällan som du vill importera sökningarna till.  
Posten <den nya datakällan> talar om att sökningarna importeras till den nya datakällan.  
Sökningar  
Här väljer du sökningarna som du vill importera till datakällan.  
Alla  
Klicka här om du vill markera alla sökningar.  
Inga  
Klicka här om du inte vill markera någon sökning.  
Till sidan Sammanfattning  
%PRODUCTNAME 5.2 databasimport - Sammanfattning  
Här ser du en sammanfattning av åtgärderna som AutoPiloten kommer att utföra.  
Dessutom kan du ge den nya datakällan ett namn.  
Ny datakälla  
Namn  
Mata in ett namn som datakällan registreras med i %PRODUCTNAME.  
Öppna den nya datakällan för administration efter importen  
Markera den här rutan om den nya datakällan ska öppnas för administration efter importen.  
Under Verktyg - Datakällor kan du administrera datakällorna.  
Adressdatakälla  
AutoPilot startar automatiskt första gången du startar %PRODUCTNAME.  
Här kan du registrera en adressbok som datakälla i %PRODUCTNAME.  
Du kan även när som helst registrera adressdata och andra datakällor i %PRODUCTNAME utan den här AutoPiloten:  
Välj typen för din externa adressbok  
Mozilla / Netscape 6.x  
Välj det här alternativet om du redan använder en adressbok i Mozilla eller Netscape 6.x.  
LDAP-adressdata  
Välj det här alternativet om du redan använder en adressbok på en LDAP-server.  
Outlook-adressbok  
Välj det här alternativet om du redan använder en adressbok i Microsoft Outlook (inte Outlook Express).  
Windowssystemets adressbok  
Välj det här alternativ om du redan använder en adressbok i Microsoft Outlook Express.  
Annan extern datakälla  
Välj det här alternativet om du vill registrera en annan datakälla som adressbok i %PRODUCTNAME nu.  
Avbryt  
Med det här kommandot avslutar du AutoPiloten utan att göra ändringar.  
Gå till föregående redigeringssteg.  
Gå till nästa redigeringssteg.  
Färdigställ  
Det här kommandot skapar anslutningen av datakällan och stänger dialogrutan.  
Ytterligare inställningar  
Här öppnar du en dialogruta där du kan göra fler inställningar.  
Inställningar  
Den här kommandoknappen öppnar en dialogruta där du kan göra fler inställningar.  
Om du har valt LDAP på den första sidan visas fliken LDAP.  
Om du har valt Annan extern datakälla på den första sidan visas en del av dialogrutan Administrera datakällor.  
Välj tabell  
Här väljer du en tabell från adressbokskällan Mozilla / Netscape 6.x som används som adressbok i %PRODUCTNAME.  
Alla tabeller från den första användarprofilen registreras för den här datakällan i %PRODUCTNAME.  
Här definierar du en av dem som den tabell som t.ex. används i fältkommandona i %PRODUCTNAME -mallarna för standardbrev (kopplad utskrift).  
Om du vill registrera tabeller från en annan användarprofil hittar du en handledning på http: / /dba.openoffice.org / howto / mozillaprofile.html.  
Listruta  
Välj ut tabellen som ska användas som adressbok i %PRODUCTNAME -mallarna.  
Det går att göra ändringar i efterhand i mallarna och dokumenten via kommandot Redigera - Byt databas.  
Datakällrubrik  
Här anger du en rubrik under vilken datakällan listas i Explorer för datakällor.  
Rubrik  
Mata in en rubrik under vilken datakällan listas i Explorer för datakällor.  
Fälttilldelning  
Här öppnar du en dialogruta där du kan definiera fälttilldelningen.  
Fälttilldelning  
Den här kommandoknappen öppnar dialogrutan Mallar: adressbokstilldelning.  
Sökningar  
Sökningar är speciella tabellvyer som t.ex. bara visar vissa poster eller några få fält per datapost och som också kan sortera dem.  
En sökning kan både gälla en tabell eller flera tabeller om de är länkade via gemensamma datafält.  
Syftet med sökningar är att enligt vissa kriterier ta fram ett särskilt urval av dataposter ur tabeller.  
Samtliga sökningar som skapats för en databas listas under databasposten Sökningar.  
Eftersom den här posten innehåller sökningar från databasen kallas den också "sökningscontainer".  
Skriva ut sökning  
För att skriva ut en sökning eller en tabell gör du så här:  
Öppna ett textdokument (eller ett tabelldokument, om du föredrar de specifika utskriftsfunktionerna för ett tabelldokument).  
Öppna databasen så att du ser sökningens namn eller tabell som post.  
Dra namnet till det öppnade dokumentet.  
Dialogrutan Infoga databaskolumner visas.  
Bestäm vilka kolumner = datafält som du vill använda.  
Klicka eventuellt på kommandoknappen AutoFormat och välj en lämplig formatering.  
Stäng dialogrutan.  
Sökningen eller tabellen infogas i dokumentet.  
Om du vill kan du göra fler ändringar och skriva ut dokumentet.  
Du kan också markera hela databastabellen i datakällvyn (kommandoknappen i hörnet av tabellen uppe till vänster) och sedan dra den till ett text - eller tabelldokument.  
I %PRODUCTNAME -hjälpen finns det mer information om att:  
Skapa ny sökning  
Om du vill skapa en ny sökning väljer du Nytt på en sökningscontainers snabbmeny.  
Sortera och filtrera data  
Om du vill ändra datavyn i en sökningstabell kan du använda sorterings - och filterfunktionerna.  
Sökningsutkast  
I fönstret Sökningsutkast kan du söka i tabeller på många olika sätt.  
Du skapar ett SQL-kommando interaktivt, som du dessutom kan redigera i efterhand.  
Sökning i flera tabeller  
Sökresultatet kan bestå av data ur flera tabeller om dessa länkats till varandra med lämpliga datafält.  
Formulera sökkriterier  
Här förklaras vilka operatorer och kommandon du kan använda när du formulerar filtervillkoren för en sökning.  
Utföra funktioner  
Du kan utföra räkneoperationer med data ur en tabell och spara resultaten som sökningsresultat.  
%PRODUCTNAME och SQL  
%PRODUCTNAME "förstår" SQL.  
Vilken syntax som ska användas beror på vilket databassystem du använder dig av.  
Element som saknas  
Där kan du välja vad som ska göras i fortsättningen.  
Hur vill du fortsätta?  
Det finns 3 alternativ för att svara på denna fråga.  
Trots detta öppna sökningen i den grafiska visningen  
Med detta alternativ öppnas sökningen i utkastvyn fastän vissa element saknas.  
När Du väljer detta alternativ kan Du dessutom ange om övriga fel ska ignoreras (se nedan).  
Sökningen öppnas i utkastvyn (det grafiska gränssnittet).  
Saknade tabeller visas tomma och ogiltiga fält visas med sitt (ogiltiga) namn i fältlistan.  
Detta ger Dig möjlighet att redigera exakt de ställen som har orsakat felet, t ex att infoga omdöpta tabeller under deras nya namn.  
Öppna sökningen i SQL-vyn  
Med det här alternativet öppnas sökningsutkastet i SQL-läge t och sökningen tolkas som Native-SQL.  
Native-SQL-läget kan först lämnas när %PRODUCTNAME kan tolka satsen fullständigt (vilket bara är möjligt om de tabeller eller fält som används i sökningen verkligen existerar).  
Öppna inte sökningen (dvs. det samma som 'Avbryt')  
Välj detta alternativ om Du vill avbryta proceduren och sökningen inte ska öppnas.  
Detta alternativ har motsvarande funktion som kommandoknappen Avbryt i dialogrutor.  
Ignorera även alla ytterligare liknande fel  
När Du har valt det första alternativet och vill öppna sökningen i den grafiska vyn trots att det saknas element, kan Du här dessutom ange om övriga fel ska ignoreras.  
Då visas inget ytterligare felmeddelande under den aktuella öppningsproceduren om sökningen inte kan tolkas korrekt.  
Sökningsutkast  
I en söknings utkastvy kan du skapa en ny sökning eller redigera en sökning som redan finns.  
Olika databaser stödjer även att en ny tabellvy skapas.  
Om du väljer Nytt vyutkast på snabbmenyn i en tabellcontainer till en sådan databas öppnas fönstret Vy, som liknar fönstret Sökning som beskrivs här.  
Utkastvyn  
När du skapar en sökning börjar du med att välja tabeller, som innehåller de data som är relevanta för sökningen.  
De här tabellerna visas i utkastvyns övre del.  
Här kan du också definiera relationer som kan förekomma mellan olika tabeller.  
Utkastvyns nedre del används för den egentliga sökningsdefinitionen.  
Här bestämmer du vilka datafält som ska användas till sökningen och efter vilka kriterier de här fälten ska visas.  
Uppe i sökningsutkastet finns det ett antal ikoner.  
Du kan t.ex. köra en skapad sökning härifrån.  
Lägg till tabeller  
När du öppnar sökningsutkastet för första gången för att skapa en ny sökning kan du klicka på Lägg till tabeller.  
En dialogruta öppnas där du kan välja de tabeller på vilka du vill basera en sökning.  
I tabellfönstret listas datafälten i de valda tabellerna.  
När du designar sökningen kan du inte ändra de tabeller som valts ut för sökningen.  
På så sätt säkerställs att tabellerna inte kan ändras när sökningen skapas.  
Även om du valt en tabell och sedan omedelbart tar bort den är den spärrad för tabellutkastet.  
Ta bort tabeller  
För att ta bort en tabell från utkastvyn klickar du på tabellfönstrets övre kant och öppnar snabbmenyn.  
Med kommandot Radera tar du bort tabellen från utkastvyn.  
Du kan också använda tangenten Delete.  
Flytta tabeller och ändra tabellstorlek  
Du kan placera tabellerna som du vill och även ändra deras storlek.  
När du ska flytta en tabell tar du tag i dess övre kant med musen och drar den till önskad position.  
För att förstora eller förminska framställningen drar du i kanten eller ett hörn.  
Relationer mellan tabeller  
Om det finns datarelationer mellan ett datafält i en tabell och ett datafält i en annan tabell kan du använda de här relationerna för din sökning.  
Om du t.ex. har en artikeltabell där varje artikel identifieras av ett entydigt artikelnummer och en kundtabell där du registrerar alla artiklar som en kund beställer och även där använder artikelnumret, finns det en relation mellan datafälten "Artikelnummer" i respektive tabell.  
Om du nu vill skapa en sökning som innehåller alla artiklar som en kund har beställt måste du hämta data ur två tabeller.  
Du talar då om för %PRODUCTNAME på vilket sätt data i den ena tabellen står i relation till data i den andra tabellen.  
Klicka på ett datafält i en tabell (t.ex. på datafältet "Artikelnummer "från kundtabellen) och dra det sedan, samtidigt som du håller ner musknappen, till datafältet i den andra tabellen ("Artikelnummer" ur artikeltabellen).  
När du nu släpper musknappen ser du en linje som förbinder de båda fälten i de båda fönstren.  
I den SQL-sökning som resulterar ur detta anges ett villkor som innebär att innehållet i båda datafälten ska var lika.  
Det går bara att skapa en sökning som baserar sig på flera tabeller som står i en relation till varandra om du använder %PRODUCTNAME som gränssnitt till en relationsdatabas, som t.ex. Adabas.  
Du kan inte söka i tabeller från olika databaser i en och samma sökning.  
Sökningar som sträcker sig över flera olika tabeller kan bara göras inom samma databassystem.  
Bestämma typ av länkning  
Om du dubbelklickar på en förbindelselinje mellan två länkade fält kan du i dialogrutan Förbindelseegenskaper bestämma typen av länkning.  
Radera relationer  
Om du vill radera en relation mellan två tabeller klickar du med musen på förbindelselinjen och trycker sedan på tangenten Delete.  
Definiera sökning  
I utkastvyns nedre del definierar Du en sökning.  
Varje kolumn i utkasttabellen innehåller ett datafält för sökningen.  
I tabellens rader kan Du för varje enskilt datafält definiera de villkor enligt vilka sökningen ska skapas.  
Villkoren på en rad knyts samman med ett logiskt OCH.  
Definiera datafält  
Markera till att börja med alla datafält i den tabell som omfattas av sökningen.  
Du kan antingen göra detta genom att dra och släppa eller genom att dubbelklicka på ett datafält i tabellfönstret.  
Att dra och släppa innebär att Du med musen drar ett datafält i ett tabellfönster till sökningsutkastets nedre del.  
Du kan bestämma i vilken kolumn respektive fält ska placeras.  
Väljer Du ett datafält genom att dubbelklicka placeras det i nästa lediga kolumn.  
Radera datafält  
Om Du vill radera ett datafält ur sökningen klickar Du med musen på fältets kolumnhuvud och ge sedan kommandot Radera i kolumnens snabbmeny.  
Spara sökning  
Du sparar sökningen med ikonen Spara på funktionslisten.  
En dialogruta öppnas där du anger ett namn för sökningen.  
Om databasen stöder scheman kan du också ange ett schema:  
Schema  
Ange namnet på schemat som tilldelas sökningsvyn / tabellvyn.  
Namn på sökning / tabellvy  
Ange namnet på sökningsvyn / tabellvyn.  
Filtrering av data  
När Du ska filtrera data för sökningen gör Du inställningar för detta i utkastvyns nedre del.  
Följande rader är tillgängliga:  
Fält  
Här anges namnet på det datafält som Du refererar till i sökningen.  
Samtliga inställningar som Du gör på de nedre raderna hänför sig till detta fält.  
När Du aktiverar en cell genom att klicka med musen visas en pilknapp med vilken Du kan välja ett fält.  
Kriteriet gäller då alla fält i tabellen.  
Alias  
Denna anges istället för ett fältnamn i en sökning.  
På så vis kan Du använda användardefinierade kolumnbeteckningar.  
Om datafältet t ex har beteckningen "ArtikelNr" och om Du istället vill att det ska visas "Artikel-nummer "i sökningen, anger Du "Artikel-nummer" som alias (utan citattecken).  
I en SQL-anvisning bestäms aliasnamn på följande sätt:  
SELECT column AS alias FROM table.  
Alltså, t ex  
SELECT "ArtikelNr" AS Artikel-Nummer FROM "Artikel "  
Tabell  
Här visas databastabellen till det valda datafältet.  
När Du aktiverar cellen genom att klicka med musen visas en pilknapp med vilken Du kan välja en annan tabell i den aktuella sökningen.  
Sortering  
Om Du klickar på cellen kan Du välja mellan sorteringsalternativen stigande, fallande eller ingen sortering alls.  
Fält av datatypen Text sorteras alfabetiskt (A till Ö) och numeriska fält sorteras numeriskt (0 till 9).  
Synlig  
Välj egenskapen Synlig för ett datafält om fältet ska synas i sökningen.  
Om du bara vill använda ett datafält för att formulera ett villkor behöver du inte visa det för sökningen.  
Kriterium  
Här anger Du ett kriterium enligt vilket innehållet i datafältet ska filtreras.  
eller  
Här kan Du ange ett kriterium för filtreringen på varje rad.  
Flera kriterier i en kolumn länkas med en ELLER-länk.  
Därutöver kan Du via radhuvudenas snabbmeny infoga en rad för funktioner i sökningsutkastets nedre del:  
Funktioner  
Här kan Du välja en funktion som ska utföras i sökningen.  
I sökningar kan Du utföra olika funktioner, beroende på vilket databassystem Du använder.  
När det gäller databaser i Adabas-format innehåller listfältet på raden Funktion följande alternativ som Du kan välja bland (aktivera visningen av raden Funktion på snabbmenyn):  
Alternativ  
SQL  
Effekt  
ingen funktion  
-  
Ingen funktion utförs  
Genomsnitt  
AVG  
Beräknar det aritmetiska medelvärdet hos ett fält.  
Antal  
COUNT  
Tomma fält räknas antingen med (a) eller inte med (b).  
a) COUNT(*):  
Om Du anger en asterisk som argument räknas alla dataposter i tabellen.  
b) COUNT(column):  
Om Du anger ett datafält som argument räknas bara de fält i vilka respektive datafält innehåller ett värde.  
Null-värden (tomma fält) räknas inte med i detta fall.  
Maximum  
MAX  
Beräknar det högsta värdet hos ett fält.  
Minimum  
MIN  
Beräknar det lägsta värdet hos ett fält.  
Summa  
SUM  
Beräknar summan av värdena hos ett fält.  
Gruppering  
GROUP BY  
Funktionerna utförs för de definierade grupperna.  
I SQL motsvarar denna inställning instruktionen GROUP BY.  
Om ett kriterium läggs till visas denna inmatning i SQL efter HAVING.  
Du kan också skriva in funktionsanrop i SQL-satsen.  
Syntaxen lyder:  
SELECT FUNCTION( column) FROM table.  
I SQL ser t ex funktionsanropet för beräkning av summa ut på följande sätt:  
SELECT SUM( "Pris") FROM "Artikel ".  
Bortsett från funktionen Gruppering rör det sig vid de ovanstående funktionerna om s.k. aggregatfunktioner.  
Det är funktioner som genom beräkningar sammanfattar data till resultat.  
Fler funktioner som inte finns med i listrutan är möjliga.  
Information om drivrutinsspecifika funktioner finns i dokumentationen till databassystemet.  
De visas sedan automatiskt på raden Funktion.  
För funktionsanrop kan Du också tilldela aliasnamn.  
Om sökningen inte ska visa funktionsnamnet i kolumnhuvudet, anger Du önskat namn under Alias.  
I en SQL-sats ser ett motsvarande funktionsanrop ut på följande sätt:  
SELECT FUNCTION() AS alias FROM table  
Exempel:  
SELECT COUNT( *) AS Antal FROM "Artikel "  
Om Du utför en funktion kan Du inte infoga ytterligare kolumner för sökningen, såvida inte dessa kolumner får funktionen "Gruppering".  
Exempel  
I följande exempel görs en sökning i två tabeller: tabellen "Artikel" med fältet "Artikel_Nr "och tabellen "Leverantörer" med fältet "Leverantör_Namn ".  
Därutöver har de båda tabellerna det gemensamma datafältet "Leverantör_Nr"  
För att kunna skapa en sökning som innehåller alla leverantörer som levererar mer än en artikel krävs följande steg:  
Infoga tabellen "Artikel" och "Leverantörer "i sökningsutkastet.  
Länka fälten "Leverantör_Nr" i båda tabellerna, såvida det inte redan finns en motsvarande relation mellan tabellerna.  
Dubbelklicka på fältet "Artikel_Nr" i tabellen "Artikel ".  
Visa raden Funktion med snabbmenyn och välj funktionen Antal.  
Ange >3 som kriterium och dölj synlig-fältet.  
Dubbelklicka på fältet "Leverantör_Namn" från tabellen "Leverantörer "och välj funktionen Gruppering.  
Utför sökningen.  
Klart!  
Om tabellen "Artikel" innehåller fälten "Pris "(pris per styck för en artikel) och "Leverantör_Nr" (för leverantörerna av artiklarna) kan Du räkna fram genomsnittspriset för artiklarna från en leverantör med följande sökning.  
Infoga tabellen "Artikel" i sökningsutkastet.  
Dubbelklicka på fälten "Pris" och "Leverantör_Nr ".  
Visa raden Funktion och välj funktionen Genomsnitt vid fältet "Pris".  
Om så önskas anges aliasnamnet "Genomsnitt" (utan citattecken) på raden för aliasnamn.  
Vid fältet "Leverantör_Nr" väljs grupperingen.  
Utför sökningen.  
Klart!  
Följande snabbmenykommandon och ikoner finns:  
Funktioner  
Visar eller döljer en rad för funktioner.  
Tabellnamn  
Visar eller döljer raden för tabellnamnet.  
Aliasnamn  
Visar eller döljer raden för aliasnamnet.  
Entydiga värden  
Om det här kommandot är aktivt överförs bara entydiga värden till sökningen.  
Av detta berörs dataposter som innehåller data som förekommer flera gånger i de valda fälten.  
I annat fall visas alla dataposter som uppfyller sökkriteriet (ALL).  
Om Du i en sökning t ex vill lista alla efternamn som förekommer i Din adressdatabas och om namnet "Svensson" förekommer flera gånger kan Du med kommandot Entydiga värden ange att namnet "Svensson "bara får förekomma en gång i sökningen.  
Vid en sökning i flera fält måste kombinationen av värden ur alla fält vara entydig för att en viss datapost ska tas med i resultatet.  
Om Du i adressboken t ex har 1x "Svensson i Stockholm" och 2x "Svensson i Göteborg "och omsökningen görs med de båda fälten "Efternamn" och "Ort "ger sökningen med kommandot Entydiga värden 1x "Svensson i Stockholm" och 1x "Svensson i Göteborg ".  
I SQL motsvarar detta kommando predikatet DISTINCT.  
Formulering av filtervillkor  
Tillsammans med jämförelseoperatorerna finns det SQL-specifika kommandon som söker innehållet i databasfält.  
När du använder de här kommandona i %PRODUCTNAME -syntax omvandlar %PRODUCTNAME dem automatiskt till motsvarande SQL-syntax.  
Du kan naturligtvis också mata in SQL-kommandot direkt.  
De följande tabellerna ger en överblick över operatorerna och kommandona:  
Operator  
Betydelse  
Villkoret är uppfyllt när...  
=  
lika med  
... fältinnehållet är identiskt med det angivna uttrycket.  
Operatorn = visas inte i sökningsfälten; om du anger ett värde utan operator används operatorn =.  
<>  
inte lika med  
... fältinnehållet inte motsvarar det angivna uttrycket.  
>  
större än  
... fältinnehållet är större än det angivna uttrycket.  
<  
mindre än  
... fältinnehållet är mindre än det angivna uttrycket.  
>=  
större än eller lika med  
... fältinnehållet är större än eller lika med det angivna uttrycket.  
<=  
mindre än eller lika med  
... fältinnehållet är mindre än eller lika med det angivna uttrycket.  
%PRODUCTNAME -kommando  
SQL-kommando  
Betydelse  
Villkoret är uppfyllt när...  
ÄR TOM  
IS NULL  
är tom  
... datafältet är tomt.  
Vid Ja / Nej-fält med tre tillstånd frågar detta kommando efter det obestämda tillståndet (varken Ja eller Nej).  
ÄR INTE TOM  
IS NOT NULL  
är inte tom  
... datafältet är inte tomt.  
SOM  
(Platshållare * för godtyckligt antal tecken  
Platshållare? för exakt ett tecken)  
LIKE  
(Platshållare% för godtyckligt antal tecken  
Platshållare _ för exakt ett tecken)  
är del av  
... datafältet innehåller det angivna uttrycket.  
Platshållare (*) anger om uttrycket x förekommer i början (x*), slutet (*x) eller inom ett fältinnehåll (*x*).  
Som platshållare kan du i SQL-sökningar ange SQL-tecknet% och i %PRODUCTNAME -gränssnittet kan du ange de platshållare du är van vid från filsystemet (*).  
Platshållaren * eller% står för ett godtyckligt antal tecken.  
För exakt ett tecken används i %PRODUCTNAME -gränssnittet frågetecknet (?) eller i SQL-sökningar understrecket (_) som platshållare.  
INTE SOM  
NOT LIKE  
är inte en del av  
... datafältet innehåller angivet uttryck.  
MELLAN x OCH y  
BETWEEN x AND y  
ligger i intervallet [x,y]  
... datafältet innehåller ett värde som ligger mellan de båda värdena x och y  
INTE MELLAN x OCH y  
NOT BETWEEN x AND y  
ligger inte i intervallet [x,y]  
... datafältet innehåller ett värde som inte ligger mellan de båda värdena x och y.  
I (a; b; c;...)  
Var noga med att semikolon används som skiljetecken i alla värdelistor.  
IN (a, b, c...)  
innehåller (a, b, c...)  
... datafältet innehåller ett av de angivna uttrycken a, b, c,...  
Sökningsresultatet fås fram med en Eller-länkning.  
Uttrycken a, b, c... kan vara siffror, men även andra tecken  
INTE I (a; b; c;...)  
NOT IN (a, b, c...)  
innehåller inte a, b, c...  
... datafältet innehåller inte ett av de angivna uttrycken a, b, c,...  
= SANN  
= TRUE  
har värdet True  
... datafältet har värdet True.  
= FALSK  
= FALSE  
har värdet False  
... datafältet har värdet False.  
Exempel  
=' Kvinna '  
returnerar datafält med fältinnehållet "Kvinna".  
SOM 'H?llo'  
returnerar datafält med fältinnehåll som "Hallo" och "Hello ".  
SOM 'S*'  
returnerar datafält med fältinnehåll som "Sun".  
MELLAN 10 OCH 20  
returnerar datafält med fältinnehåll med värden mellan 10 och 20. (Det kan både röra sig om textfält och sifferfält).  
I (1; 3; 5; 7)  
returnerar datafält med värdena 1, 3, 5, 7.  
Innehåller datafältet t.ex. ett artikelnummer kan du skapa en sökning som tar fram vissa artiklar med det angivna numret.  
INTE I ('Svensson')  
returnerar datafält som inte innehåller "Svensson".  
Datumfält visas generellt i formatet #Datum# så att de entydigt ska kunna identifieras som datum.  
Datumvillkoret avbildas på följande ODBC-kompatibla sätt i den resulterande SQL-satsen.  
Datum  
{D'YYYY-MM-DD'}  
Datumtid  
{D'YYYY-MM-DD HH:MM:SS'}  
Tid  
{D'HH:MM:SS'}  
Dessutom stöder %PRODUCTNAME följande Escape-sekvenser som förekommer i ODBC och JDBC.  
Datum  
{d 'YYYY-MM-DD'}  
Tid  
{t 'HH:MI:SS[.SS]'} - [] optional  
Datumtid  
{ts 'YYYY-MM-DD HH:MI:SS[.SS]'} - [] optional  
Exempel: select {d '1999-12-31'} from world.years  
Like Escape Sequence: {escape 'escape-character'}  
Exempel: select * from Artikel where Artikelnamn like 'The *%' {escape '*'}  
Exemplet ger alla poster där artikelnamnet börjar med "The *".  
På så sätt kan Du också söka efter tecken som i vanliga fall tolkas som platshållare, t ex *,?, _,% eller punkt.  
Outer Join Escape Sequence: {oj outer-join}  
Exempel: select Artikel.* from {oj Artikel LEFT OUTER JOIN Beställningar ON Artikel.Nr=Beställningar.ANR}  
I annat fall utvärderas de som en teckenföljd (sträng). 'Strängar 'omges av enkla citattecken.  
Sökning i textfält  
För att söka innehållet i ett textfält ska uttrycket sättas inom enkla citattecken.  
Det görs ingen åtskillnad mellan versaler och gemener.  
Sökning i datumfält  
Även när Du vill filtrera fram ett visst datum anger Du uttrycket inom enkla citattecken.  
Följande format kan användas:  
ÅÅÅÅ-MM-DD TT:MM:SS och ÅÅÅÅ / MM / DD TT:MM:SS liksom även ÅÅÅÅ.MM.DD TT:MM:SS  
Sökningar i Ja / Nej-fält  
För att göra sökningar i Ja / Nej-fält använder Du vid dBase - eller Adabas - tabeller följande syntax:  
Tillstånd  
Sökningskriterium  
Exempel  
Ja  
för dBase-tabeller: ett godtyckligt värde ej lika med 0  
=1 ger alla dataposter för vilka Ja / Nej-fältet har tillståndet "Ja" eller "Till "(svart markering)  
Nej  
0  
=0 ger alla dataposter för vilka Ja / Nej-fältet har tillståndet "Nej" eller "Från "(ingen markering)  
Tom  
IS NULL respektive ÄR TOM  
IS NULL ger alla dataposter för vilka Ja / Nej-fältet inte intar något av tillstånden Ja eller Nej (grå markering).  
Vilken syntax som ska användas beror på vilket databassystem Du använder.  
Tänk också på att Ja / Nej-fält kan vara definierade på olika sätt (inte 3, utan 2 tillstånd).  
Parametersökningar  
Alternativt kan Du använda ett likhetstecken med kolon (=:x).  
När sökningen utförs får Du i en dialogruta en fråga om vilket uttryck variabeln x ska tilldelas.  
Om Du söker efter parametrar visas i dialogrutan en listruta med alla parametrar och bredvid varje parameter en inmatningsrad.  
Det bästa sättet är att ange värdena uppifrån och ned och att efter varje värde trycka på returtangenten.  
Det går inte att göra parametersökningar med platshållare (*,_) eller specialtecken (?, o.s.v.)  
Om du vill formulera en parametersökning och spara den med variablerna kan du senare lätt skapa en sökning där du bara behöver ersätta variablerna med de önskade uttrycken. %PRODUCTNAME frågar efter de här variablerna i en dialogruta, så snart du öppnat sökningen.  
Ange parametervärde  
I denna dialogruta söks de variabler som Du definierat i sökningen.  
Bekräfta inmatningen med OK.  
Parametersökningar krävs också för underformulär, eftersom dessa uteslutande arbetar med sökningar vid vilka de värden som hämtas internt läses ur en variabel.  
I SQL-satsen ser en parametersökning t.ex. ut så här:  
select * from 'adressen' where 'name '= :placeholder  
SQL-läge  
SQL står för "Structured Query Language" och är ett språk som används för att ställa frågor till, uppdatera och hantera relationsdatabaser.  
I %PRODUCTNAME behöver du sällan SQL-kunskaper när du gör sökningar, eftersom du inte behöver ange någon SQL-kod.  
När du skapar en sökning i sökningsutkastet omvandlar %PRODUCTNAME automatiskt dina anvisningar till motsvarande SQL-syntax.  
Om du byter SQL-vy du med hjälp av ikonen Sätt på / stäng av designvy kan du se SQL-kommandona för en sökning som har skapats.  
Du kan formulera din sökning direkt i SQL-kod.  
Men tänk på att den speciella syntaxen beror på vilket databassystem du använder.  
Adabas-formatet baserar sig på standarden SQL / 92 (ofta kallad SQL2), som lanserades 1989 av ISO och flera nationella standardiseringsorganisationer (särskilt ANSI) och utvidgades 1992.  
Om du matar in SQL-koden manuellt kan du skapa SQL-specifika sökningar som inte stöds av det grafiska gränssnittet i Sökningsutkast et.  
De här sökningarna måste i göras i Native-SQL-läge.  
Genom att klicka på ikonen Utför SQL-kommando direkt i SQL-vyn kan du formulera en sökning som inte bearbetas av %PRODUCTNAME.  
För databaser i Adabas-format gäller följande konventioner för SQL-syntax:  
Tabell - och kolumnnamn sätts inom dubbla citattecken och strängar identifieras av enkla citattecken.  
Aliasnamn ges ingen speciell markering.  
Egenskaper för sammanslagning (join)  
Om du dubbelklickar på en förbindelselinje mellan två länkade fält i sökningsutkastet, kan du definiera typ av länk i dialogrutan Egenskaper för sammanslagning (join).  
Den här inställningen används sedan för alla sökningar som skapas.  
Alternativ  
Här kan du definiera av vilken typ den valda sammanslagningen ska vara.  
Det som skiljer sökningar med de olika länkningstyperna är antalet dataposter som visas.  
Du kan välja mellan fyra alternativ:  
Inre  
Vid inre join innehåller resultattabellen bara de dataposter där innehållet i de länkade fälten är lika.  
I SQL i %PRODUCTNAME åstadkoms denna jointyp genom en motsvarande WHERE-instruktion.  
Vänster  
Vid vänster join innehåller resultattabellen alla fält ur den vänstra tabellen och ur den högra tabellen bara de fält hos vilka innehållet i de länkade fälten är lika.  
I SQL i %PRODUCTNAME motsvarar den här jointypen kommandot LEFT OUTER JOIN.  
Höger  
Vid höger join innehåller resultattabellen alla fält ur den högra tabellen och ur den vänstra tabellen bara de fält hos vilka innehållet i de länkade fälten är lika.  
I SQL i %PRODUCTNAME motsvarar den här jointypen kommandot RIGHT OUTER JOIN.  
Fullständig  
Vid fullständig join innehåller resultattabellen alla fält ur den vänstra och den högra tabellen.  
I SQL i %PRODUCTNAME motsvarar den här jointypen kommandot FULL OUTER JOIN.  
Visningsfält  
Visar hjälp till det valda alternativet.  
Formulär  
Formulär använder du för att komma åt data i en tabell, och du kan använda dem till att lägga in nya data eller ändra befintliga data.  
Till skillnad mot datavyn i en tabell, visar ett formulär bara en datapost åt gången och bara de fält som du har valt.  
Samtliga formulär som har skapats till en databas med %PRODUCTNAME listas under databasposten Formulär.  
Eftersom den här posten innehåller databasens formulär kallas den också "formulärcontainer".  
Formulär som du skapar i ett %PRODUCTNAME -dokument med hjälp av kommandona på utrullningslisten Formulär kan du spara var som helst som vanliga dokument.  
De här formulären visas inte i formulärcontainern i %PRODUCTNAME, utan behandlas som dokument av respektive typ.  
I %PRODUCTNAME -hjälpen finns det mer information om att:  
Skapa ett nytt formulär  
Om du vill skapa ett nytt formulär väljer du Nytt på formulärcontainerns snabbmeny.  
AutoPilot  
Här hittar du en noggrann beskrivning av de sidor i AutoPiloten som visas när du skapar ett formulär.  
Formulärfunktioner  
Formulärfunktionerna ger dig alla verktyg som du behöver för att skapa ett formulär i ett text-, tabell-, tecknings - eller presentationsdokument.  
Formulär i utkastläge  
I utkastläget skapar du ett formulär och definierar framför allt formulärets egenskaper och kontrollfälten som det innehåller.  
Sortera och filtrera data  
Sorterings - och filterfunktionerna hittar du på formulärlisten när du har öppnat ett formulär i användarläge.  
Underordnat formulär  
Snabbmenyer till formulär  
På formulärcontainerns snabbmeny finns olika funktioner som gäller allmänt för alla formulär i databasen.  
Om du vill redigera ett speciellt formulär i databasen, markerar du det och öppnar sedan den tillhörande snabbmenyn.  
På snabbmenyerna hittar du följande kommandon:  
Nytt  
Om ett formulär är markerat kommer du till formulärvyn.  
På snabbmenyn till ett speciellt formulär visas dessutom följande kommandon:  
Formulärutkast  
Detta kommando öppnar formuläret i utkastläge.  
För skrivskyddade databaser är detta kommando inte tillgängligt.  
Formulär raderas fysiskt.  
Nytt formulär  
Välj Nytt formulär på en "Länkar "-post i Explorer för datakällor om du vill skapa ett nytt formulär.  
Då öppnas en undermeny där du kan välja om du vill skapa formuläret med hjälp av en AutoPilot eller om det ska skapas i ett text-, tabell - eller presentationsdokument.  
Om du väljer ett av kommandona Textdokument, Tabelldokument eller Presentation, måste du skapa formuläret manuellt.  
Ett tomt dokument av respektive typ öppnas där du kan använda formulärfunktionerna för att utforma formuläret i den önskade miljön.  
Om du väljer Från mall visas sedan dialogrutan Mallar och dokument där du kan välja en mall som används som utgångspunkt för formuläret.  
Infoga de önskade formulärfunktionerna och spara det nya formuläret.  
Om du väljer AutoPilot, guidas du sedan av en assistent genom de olika stegen för att skapa ett nytt formulär.  
Spara formulär  
Här anger du med vilket namn objektet ska sparas.  
När du klickar på OK visas det nya objektet med sitt namn i databasens motsvarande container.  
Om du skapar ett formulär i ett text-, tabell - eller presentationsdokument, öppnas dialogrutan Spara som när du sparar dokumentet första gången.  
Här anger du med vilket namn formuläret ska sparas.  
När du klickar på OK visas en motsvarande post för det nya formuläret i databasens formulärcontainer.  
Om du använder AutoPiloten för att skapa ett nytt formulär, så sparas formuläret så snart du klickar på kommandoknappen Färdigställ på assistentens sista sida.  
Formuläret visas sedan också under sitt namn i datakällans "Länkar "-container.  
Formulärutkast  
Alla %PRODUCTNAME -dokument kan göras till ett formulär.  
Foga bara in en eller flera formulärfunktioner.  
På verktygslisten finns ikonen Formulär.  
Den öppnar en utrullningslist med samtliga grundläggande funktioner som behövs för redigering av formuläret.  
Många av de här funktionerna hittar du även på objektlisten om du markerar ett formulärelement.  
När du klickar på ett formulärelement i redigeringsläget får du tillgång till sammanhangsanpassade redigeringsfunktioner på objektlisten, Format -menyn och snabbmenyerna.  
I formulärutkastet kan du integrera kontrollfält, tilldela dem egenskaper, definiera formuläregenskaper och definiera underordnade formulär.  
Formulär-Navigator som du öppnar via objektlisten eller utrullningslisten är ett användbart hjälpmedel.  
Med kommandot Öppna i utkastläge kan du spara ett formulärdokument på ett sådant sätt att det alltid öppnas i redigeringsläge.  
Om det uppstår ett fel när egenskaperna för de objekt som finns i formuläret ska tilldelas (t.ex. om en icke-existerande databastabell tilldelas ett objekt), så visas ett motsvarande felmeddelande.  
I detta felmeddelande kan det finnas en kommandoknapp som heter Fler.  
Nu öppnas en dialogruta som på ett översiktligt sätt visar information, varningar och fel till det aktuella problemet.  
Tabeller  
I datakällornas tabeller visas data rad för rad.  
Du kan ange data på nytt och radera data.  
I %PRODUCTNAME -hjälpen hittar du mer information om att:  
Skapa nytt tabellutkast eller redigera tabellutkast  
Sortera och filtrera data  
Relationer, primärnycklar och sekundärnycklar  
Snabbmenyer till tabeller  
På tabellcontainerns snabbmeny finns olika funktioner som gäller allmänt för alla tabeller i databasen.  
Om du vill redigera en speciell tabell i databasen, markerar du den och öppnar sedan den tillhörande snabbmenyn.  
Allt efter sammanhang kan det hända att du inte kommer att hitta alla de funktioner som nämns här för din aktuella databas.  
Kommandot Relationer, som används för att definiera relationer mellan olika tabeller, är exempelvis bara tillgängligt för relationsdatabaser.  
På snabbmenyerna hittar du, beroende på vilket databassystem som används, följande poster:  
När du har öppnat en tabell, har du tillgång till olika funktioner för att redigera data.  
Användarinställningar  
I den här dialogrutan gör du användarinställningar för en Adabas-tabell.  
Användarurval  
Här väljer du användare, lägger till eller raderar användare och ändrar lösenord.  
Användare  
Markera den användare vars inställningar du vill redigera.  
Lägg till användare  
Klicka här om du vill skapa en ny användare.  
Ändra lösenord...  
Klicka här om du vill ändra lösenordet för den markerade användaren.  
Radera användare...  
Klicka här om du vill radera den markerade användaren.  
Åtkomsträttigheter för markerad användare  
Här kan du se och tilldela rättigheter för en markerad användare.  
Mata in / ändra lösenord  
I den här dialogrutan skriver du in ett lösenord och bekräftar det.  
Om du skapar en ny användare anger du dennes namn i den här dialogrutan.  
Användare  
Här anger du namnet för den nya användaren.  
Det här fältet visas bara när du skapar en ny användare.  
Gammalt lösenord  
Här anger du det gamla lösenordet.  
Det här fältet visas om du har öppnat dialogrutan via Ändra lösenord.  
Lösenord  
Här anger du lösenordet.  
Bekräfta (lösenord)  
Här upprepar du lösenordet.  
Tabellutkast  
I Tabellutkast -fönstret definierar du nya tabeller eller redigerar en tabells struktur.  
Fönstret har en egen menylist och en egen funktionslist.  
Där finns följande nya kommando:  
Indexutkast  
Tabelldefinitionsområde  
Här definierar du tabellstrukturen.  
Fältnamn  
Ange namnet för datafältet.  
Håll dig till databasens restriktioner, t.ex. när det gäller längden på namnet, specialtecken och blanksteg.  
Fälttyp  
Välj en fälttyp.  
Beskrivning  
Ange en beskrivning om du vill.  
Snabbmenyn på radhuvudena innehåller följande kommandon:  
Klipp ut  
Klipper ut den markerade raden / de markerade raderna och placerar den / dem i urklippet.  
Kopiera  
Kopierar den markerade raden / de markerade raderna till urklippet.  
Klistra in  
Klistrar in urklippets innehåll.  
Radera  
Raderar den markerade raden / de markerade raderna.  
Infoga rader  
Så många rader som du har markerat infogas framför de markerade raderna.  
Primärnyckel  
Om det finns en bock framför kommandot är datafältet på den här raden en primärnyckel.  
Genom att klicka på kommandot aktiverar och deaktiverar du denna status.  
Kommandot visas bara om datakälan understöder primärnycklar.  
Fältegenskaper  
Här definierar du fältegenskaperna för det fält som just är markerat.  
Längd  
Ange datafältets längd.  
Antal decimaler  
Ange antalet decimaler för ett talfält eller decimalfält.  
Standardvärde  
Ange ett värde som är förinställt i nya dataposter.  
Formatexempel  
Här ser du formatbeskrivningen som du kan välja ut med hjälp av kommandoknappen....  
...  
Den här kommandoknappen öppnar dialogrutan Fältformatering.  
Hjälpområde  
Här visas hjälptexter.  
Indexutkast  
I dialogrutan Indexutkast redigerar du index för den aktuella tabellen.  
Indexlista  
I listan väljer du ett index som du vill redigera.  
Till höger i dialogrutan visas då de tillhörande indexdetaljerna.  
Nytt index  
Här skapar du ett nytt index.  
Radera aktuellt index  
Raderar det aktuella indexet.  
Byt namn på aktuellt index  
Om du klickar här kan du byta namn på det aktuella indexet i listan.  
Spara aktuellt index  
Sparar det aktuella indexet i datakällan.  
Återställ aktuellt index  
Återställer det aktuella indexets inställning som det hade när dialogrutan öppnades.  
Indexdetaljer  
När du ändrar en detalj för det aktuella indexet och sedan markerar ett annat index överförs den här ändringen direkt till datakällan.  
Du kan bara lämna dialogrutan eller markera ett annat index om ändringen har kvitterats av datakällan.  
Men du kan ångra ändringen genom att klicka på Återställ aktuellt index.  
Entydigt  
Markera den här rutan om indexet ska vara entydigt.  
Då får inga dataposter i det här datafältet ha samma innehåll.  
Fält  
Här väljer du det datafält som ska bli ett indexfält.  
Du kan också välja flera fält.  
Om du vill avmarkera ett fält väljer du den tomma posten i början av listan.  
Indexfält  
Välj ett eller flera fält.  
Sorteringsordning  
Välj sorteringsordning.  
Stäng  
Här stänger du dialogrutan.  
Du tillfrågas om du vill spara ändringarna eller inte.  
Relationer  
Det här kommandot öppnar ett fönster där du kan definiera länkar mellan olika databastabeller.  
Här kan du koppla samman tabellerna i den aktuella databasens via gemensamma datafält.  
Den här funktion är bara tillgänglig för relationsdatabassystem, d.v.s. kommandot är bara synligt om du använder %PRODUCTNAME som frontend för en relationsdatabas.  
Om du väljer Relationsutkast i tabellcontainerns snabbmeny, öppnas ett fönster där alla befintliga relationer mellan tabellerna i den aktuella databasen.  
Om det ännu inte har definierats några relationer eller om du vill sammankoppla fler tabeller i databasen, så klickar du på ikonen Lägg till tabeller.  
Sedan öppnas en dialogruta där du kan välja de önskade tabellerna.  
När relationsfönstret är öppet kan de valda tabellerna inte redigeras i tabellutkastläget.  
På så vis garanteras att tabellerna inte kan ändras i just det ögonblick då relationerna skapas.  
De valda tabellerna visas i det övre området i utkastvyn.  
Ett tabellfönster kan du ta bort igen via snabbmenyn eller med Delete-tangenten.  
Primärnyckel och sekundärnyckel  
Om du vill kunna skapa en relation mellan olika tabeller, måste det finnas minst en primärnyckel som entydigt kännetecknar ett datafält i respektive tabell.  
Då kan du från andra tabeller hänvisa till denna primärnyckel för att få åtkomst till data i den här tabellen.  
De datafält som motsvarar primärnyckeln och som hänvisar till den kallas sekundärnycklar.  
Datafält till vilka en primärnyckel har tilldelats markeras i tabellfönstret genom en liten nyckelsymbol.  
Titta exempelvis på tabellen "Artikel", där man via ett artikelnummer kan identifiera varje enskild datapost.  
Fältet "Artikelnummer" är i denna tabell alltså en entydig nyckel, en så kallad primärnyckel.  
I databasen finns det ytterligare en tabell som kallas "Beställningar".  
Till varje datapost i denna tabell tillordnas via ett fält "Artikelnummer" den beställda artikelns nummer.  
Även detta fält är ett nyckelfält.  
Det innehåller nämligen en nyckel för att få åtkomst till dataposterna i en annan tabell, i detta fall till dem i tabellen "Artikel".  
Detta fält kallas därför även för sekundärnyckel.  
Med en relation skapas en relation mellan primärnyckeln för tabellen "Artikel" och sekundärnyckeln för tabellen "Beställningar ".  
Definiera relationer  
Alla befintliga relationer visas i relationsfönstret med en linje, med vilken primär - och sekundärnyckelfälten kopplas samman.  
Du lägger till en relation genom att dra ett fält i en tabell med musen och släppa det på fältet i den andra tabellen.  
En relation tas bort igen om du trycker på Delete-tangenten (relationen måste vara markerad).  
Du kan även klicka på ikonen Ny relation i relationsfönstrets övre del och definiera relationen mellan två tabeller i en dialogruta.  
Om du använder %PRODUCTNAME som frontend för en relationsdatabas, så sparar %PRODUCTNAME inte processerna temporärt när du skapar och raderar relationer utan processerna vidarebefordras direkt till den externa databasen!  
Om du dubbelklickar på en förbindelselinje kan du tilldela relationen vissa egenskaper.  
Nu öppnas dialogrutan Relationer.  
Relationer  
Här definierar du en relation mellan två tabeller.  
De här uppdaterings - och raderingsalternativen är bara tillgängliga om de stöds av den databas som används.  
Tabeller  
Här visas de två tabeller mellan vilka det finns en relation.  
När du skapar en ny relation kan du välja vardera en tabell ur de två kombinationsfälten i den övre delen av dialogrutan.  
Om du har öppnat dialogrutan Relationer till en redan befintlig relation genom att dubbelklicka på förbindelselinjen i relationsfönstret, så kan de tabeller som ingår i relationen inte förändras här.  
Nyckelfält  
Här definierar du nyckelfält för relationen.  
Namnen på de tabeller som valts för relationen visas här som kolumnnamn.  
Om du klickar i ett fält, så kan du med hjälp av pilknappen välja ett fält i tabellen.  
Varje relation skrivs på en rad.  
Uppdateringsalternativ  
Här gör du inställningar som ska gälla när ett primärnyckelfält ändras.  
Ingen åtgärd  
Ifall detta alternativ är aktiverat och en primärnyckel ändras, påverkas inte andra sekundärnyckel-fält.  
Uppdatera kaskad  
Med detta alternativ uppdateras alla sekundärnyckel-fält om värdet för det tillhörande primärnyckel-fältet ändras (Cascading Update).  
Sätt null  
Med det här alternativet tilldelar du sekundärnyckelfälten värdet "IS NULL" om den tillhörande primärnyckeln ändras.  
IS NULL betyder här att datafältet är tomt.  
Sätt standard  
Med det här alternativet tilldelar du sekundärnyckelfälten ett standardvärde om den tillhörande primärnyckeln ändras.  
Detta standardvärde för ett sekundärnyckel-fält definierades när den tillhörande tabellen skapades och fältegenskaperna bestämdes.  
Raderingsalternativ  
Här väljer du de alternativ som ska gälla när ett primärnyckelfält raderas.  
Ingen åtgärd  
Ifall detta alternativ är aktiverat och en primärnyckel raderas, påverkas inte andra sekundärnyckel-fält.  
Radera kaskad  
Med detta alternativ raderas alla sekundärnyckel-fält om det tillhörande primärnyckel-fältet raderas (Cascading Delete).  
När det gäller detta alternativ bör du tänka på följande: när ett primärnyckelfält raderas, så raderas även alla dataposter i andra tabeller som har denna nyckel som sekundärnyckel.  
Var därför försiktig när du använder det här alternativet eftersom det i värsta fall kan leda till att en stor del av hela databasen raderas!  
Sätt null  
Med detta alternativ tilldelas sekundärnyckel-fälten värdet "IS NULL" om den tillhörande primärnyckeln raderas.  
Sätt standard  
Med detta alternativ tilldelas sekundärnyckel-fälten ett standardvärde om den tillhörande primärnyckeln raderas.  
Kopiera sökning eller tabell med dra-och-släpp  
I den här dialogrutan anger du alternativen för kopiering av en sökning eller tabell.  
Du kan kopiera en sökning från %PRODUCTNAME genom att dra och släppa, men även en tabell från ett %PRODUCTNAME Writer - eller HTML-dokument eller en markerad del av det, eller ett cellområde från en %PRODUCTNAME Calc-tabell.  
Du redigerar sökningen genom att dra och släppa.  
På så vis kan du:  
skapa en kopia av sökningen,  
överföra sökningens data till en annan sökning,  
använda tabellstrukturen som bas för en ny tabell.  
Det spelar ingen roll om utbytet ska ske inom samma databas eller mellan olika databaser.  
Markera sökningen med musen och dra den till den önskade databasens tabellcontainer.  
Kopiera tabell  
Om du kopierar en sökning eller tabell till en tabellcontainer med dra-och-släpp i datakällvyn, visas AutoPilot Kopiera tabell.  
Tabellnamn  
Här skriver du det namn med vilket kopian av objektet ska sparas på den plats du väljer.  
En del databasformat stöder bara namn med 8 tecken.  
Alternativ  
Definition och data  
Med det här alternativet skapar du en 1:1-kopia av databastabellen.  
Både tabelldefinitionen och samtliga data kopieras.  
Tabelldefinitionen omfattar tabellens struktur och uppbyggnad av olika datafält inklusive de speciella fältegenskaperna.  
Fältinnehållet bestämmer dessa data.  
Definition  
Med det här alternativet kopierar du bara tabelldefinitionen, data överförs inte.  
Som tabellvy  
Det här alternativet kan du bara välja när en sökning kopieras till en tabellcontainer, och om databasen stöder vyer (views).  
Genom det här alternativet kan du visa och redigera en sökning i en "normal" tabellvy.  
Tabellen filtreras i vyn genom SQL-satsen "Select".  
Tillfoga data  
Om du väljer det här alternativet, infogas data från den tabell som ska kopieras i en redan existerande tabell.  
En förutsättning för att den här åtgärden ska kunna genomföras med lyckat resultat är att tabelldefinitionen är identisk med de data som ska kopieras.  
Data kan inte importeras om måltabellen inte innehåller ett motsvarande datafält av samma typ.  
Du tilldelar datafältnamn på sidan Tilldela kolumner i AutoPiloten Kopiera tabell.  
Om data inte kan tillfogas helt eller delvis, visas en lista med de fält vars data inte kan importeras i dialogrutan Kolumninformation.  
Om du bekräftar den här dialogrutan genom att klicka på OK, tillfogas bara de data som uppfyller kriterierna för en lyckad kopiering.  
Om fältlängden i måltabellen är mindre än den i källtabellen, när data tillfogas, anpassas fältinnehållet i den kopierade tabellen till fältlängden i måltabellen.  
Skapa primärnyckel  
Om du markerar den här rutan skapas automatiskt ett primärnyckelfält som fylls med värden.  
Det här fältet bör du använda när du t.ex. kopierar en dBase-tabell till Adabas-format, då det alltid måste finnas en primärnyckel i Adabas-format när en tabell redigeras.  
Namn:  
Här kan du ge den skapade primärnyckeln ett namn.  
Till sidan 2 i AutoPiloten  
Överta kolumner  
Om du kopierar en sökning eller tabell med dra-och-släpp till en tabellcontainer i datakällvyn visas Autopilot Kopiera tabell.  
Detta är sidan 2 i AutoPiloten.  
Existerande kolumner  
Vänstra fältet  
I det vänstra fältet väljer du datafälten som du vill använda i måltabellen eller målsökningen.  
Klicka på >.  
Högra fältet  
Här visas datafälten som har överförts.  
Kommandoknappar  
Med > överför du fälten som har markerats på den vänstra sidan till den högra, med < överför du de fält som har markerats på den högra sidan till den vänstra.  
Med >> och << överför du alla fält.  
Till sidan 3 i AutoPiloten  
Typformateringar  
Detta är sidan 3 i AutoPiloten.  
Listruta  
Här väljer du ett datafält som du vill se kolumninformation till eller redigera.  
Kolumninformation  
Här tittar du på eller redigerar kolumninformation till ett datafält.  
Beroende på den valda fälttypen visas olika inmatningsfält.  
Fältnamn  
Här anger du namnet som datafältet ska få i den nya tabellen.  
Observera eventuella restriktioner som databasen har.  
Fälttyp  
Välj fälttyp.  
Längd  
Ange längden på datafältet.  
Antal decimaler  
Anger antalet decimaler för ett talfält eller decimalfält.  
Standardvärde  
Välj det förinställda värdet för ett Ja / Nej-fält.  
Automatisk typigenkänning  
Det här området visas om du t.ex. drar en tabell från ett dokument med dra-och-släpp till en tabellcontainer.  
Datafälttyperna kan ofta kännas igen automatiskt på innehållet.  
(max) rader  
Här anger du hur många rader som används för att uppnå en automatisk typigenkänning.  
Auto  
Med den här kommandoknappen startar du den automatiska typigenkänningen.  
Tilldela kolumner  
På den här sidan definierar du vilket datafältinnehåll i en källtabell som ska kopieras till vilka andra datafält i måltabellen.  
Dialogrutan visas som andra sida i AutoPiloten Kopiera tabell vid dra-och-släpp av tabeller när du har valt alternativet Tillfoga data på den första sidan.  
Flytta posterna på den vänstra eller högra sidan fram och tillbaka med hjälp av kommandoknapparna, tills de korresponderande datafältnamnen ligger bredvid varandra i båda listorna.  
Datafältens ordning i måltabellen ändras inte: i den här dialogrutan gäller det bara tilldelningen vid kopiering.  
Källtabell  
Här ser du alla tillgängliga datafält i källtabellen där de data som ska tillfogas kommer ifrån.  
Du kan markera datafälten vars innehåll ska kopieras i rutorna framför datafältnamnen.  
Med kommandoknapparna alla och inga kan du markera resp. avmarkera alla datafältnamn samtdigt.  
Måltabell  
Här visas alla datafält i måltabellen där nya data ska infogas.  
upp  
Den markerade posten på den här sidan i dialogrutan flyttas tillsammans med sin markering ett steg uppåt.  
På den andra sidan i dialogrutan flyttas bara markeringen, inte den markerade posten.  
ned  
Den markerade posten på den här sidan i dialogrutan flyttas tillsammans med sin markering ett steg nedåt.  
På den andra sidan i dialogrutan flyttas bara markeringen, inte den markerade posten.  
alla  
Alla poster i källtabellen får en markering.  
Allt innehåll i de markerade datafälten tillfogas måltabellen.  
inga  
Alla markeringar i källtabellen tas bort.  
Allmänt  
I egenskapsdialogrutan till en databastabell kan du bl.a. definiera de rättigheter som den aktuella användaren har för tabellen.  
Allmänt  
Om du skapar en databastabell som administratör, kan du se under den här fliken om och i vilken omfattning en användare, som har åtkomst till den här tabellen, får ändra data eller tabellstrukturen.  
Du kommer till fliken via en tabells snabbmeny - menykommandot Egenskaper.  
Som aktuell användare kan du se vilka rättigheter du har för tabellen i egenskapsdialogrutan under fliken Allmänt.  
Om du exempelvis inte får radera data i en tabell kan du se information om detta under fliken Allmänt.  
De olika egenskaperna kan du inte ändra här.  
Namn  
Här skrivs databastabellens namn in.  
Typ  
Här anges objektets typ, d.v.s. "Tabell" för databastabeller.  
Placering  
Här återges hela sökvägen för databastabellen.  
Läs data  
Om denna kryssruta är markerad, får data läsas av användaren.  
Infoga data  
Om denna kryssruta är markerad, får nya data infogas av användaren.  
Ändra data  
Om denna kryssruta är markerad, får data ändras av användaren.  
Radera data  
Om denna kryssruta är markerad, får data raderas av användaren.  
Ändra tabellstruktur  
Om denna kryssruta är markerad, får tabellstrukturen ändras av användaren.  
Radera tabellstruktur  
Om denna kryssruta är markerad, får tabellstrukturen raderas av användaren.  
Ändra referens  
Om denna kryssruta är markerad, får angivna referenser ändras av användaren.  
Det innebär att användaren får ange relationer för dessa tabeller eller radera redan existerande.  
Beskrivning  
Här visas beskrivningen som angetts för den här tabellen.  
Tabellbeskrivning  
I det här fältet visas beskrivningen för den aktuella tabellen..  
Databaser  
Du registrerar databaser som du vill använda i %PRODUCTNAME med Verktyg - Datakällor.  
Datakällor i %PRODUCTNAME  
Datakällegenskaper  
Kopiera eller flytta databasobjekt med dra-och-släpp  
Mata in SQL-kommando  
Databassystem som stöds  
Se även ytterligare information om %PRODUCTNAME -datakällor.  
Datakällor i %PRODUCTNAME  
Här finns information om hur du arbetar med datakällor i %PRODUCTNAME.  
Övrigt innehåll på denna sida:  
Adressboken  
Ställa in datakälla  
Öppna datakälla  
Kopiera eller flytta databasobjekt med dra-och-släpp  
Adressboken  
I en dialogruta kan du definiera vilket datafält från din systemadressbok som ska tilldelas vilken platshållare.  
Du kan öppna den här dialogrutan via Arkiv - Dokumentmall - Adressbokskälla; den startas dessutom automatiskt när du använder en av dokumentmallarna för första gången och den här tilldelningen inte har gjorts ännu.  
Ställa in en ny datakälla  
I en dialogruta under Verktyg - Datakällor kan du specificera datakällan och ge den ett namn med vilket den anropas i %PRODUCTNAME.  
Beroende på vald typ kan du ange olika alternativ.  
När du ställer in en befintlig databas i %PRODUCTNAME anger du helt enkelt datakällan.  
För en text - eller dBase-databas är det en mapp som innehåller databasen med dess tabeller.  
Här bildar alla tabeller (databasfiler) i en mapp (katalog) tillsammans en databas.  
När du registrerar en datakälla i %PRODUCTNAME skapas i princip bara en länk till databestånden.  
Den här länken ger dig åtkomst till data.  
Så här öppnar du en datakälla  
Datenkällvyn visas och döljs när du trycker på F4 när ett text-, tabell - eller formeldokument är öppet.  
Om du öppnar en datakälla genom att klicka på plustecknet framför datakällans namn visas posterna för länkar, sökningar och tabeller.  
Kopiera eller flytta databasobjekt med dra-och-släpp  
Internt i %PRODUCTNAME kan du flytta databasinnehåll mellan olika databaser genom att dra och släppa det med musen.  
Även inom en databas kan du lätt skapa kopior till ett databasobjekt genom att dra och släppa.  
När du exempelvis vill skapa en ny sökning som bara skiljer sig något från en redan existerande, så kan du helt enkelt kopiera denna sökning och sedan göra ändringarna i sökningsutkastet.  
Dessutom kan du dra en tabell eller markerade delar av tabeller ur ett %PRODUCTNAME Writer-dokument, ett HTML-dokument eller ur %PRODUCTNAME Calc och släppa den på en tabellcontainer.  
Det går lika bra att t.ex. dra en tabell från datakällvyn till ett textdokument.  
Databasobjekt kan du både kopiera och flytta.  
Vid kopiering bibehålls originalet, vid flyttning raderas originalet.  
Om du vill kopiera ett objekt, behöver du bara dra det med musen till det önskade stället.  
Om du vill flytta objektet, håller du samtidigt ner skifttangenten.  
Om du vill kopiera eller flytta flera databasobjekt av en typ, så markerar du dem efter varandra innan du drar dem med musen till destinationsorten.  
Vid konverteringar mellan olika databastyper måste man ta hänsyn till att fältdefinitionerna motsvarar olika konventioner.  
Fält - resp. kolumnnamn för dBase-tabeller får exempelvis bara vara 10 tecken långa, för Adabas-tabeller däremot 18.  
Om du kopierar eller flyttar en tabell genom att dra och släppa den, och om den tillåtna teckenlängden för ett fält i måltabellen är mindre än i källtabellen, så uppmanas du i en dialogruta att ange ett nytt fältnamn.  
Du kan även använda Auto-knappen i den här dialogrutan, då anpassas namnen automatiskt av %PRODUCTNAME.  
Kopiera eller flytta sökning  
Om du drar och släpper en sökning, så kopieras sökningen om du släpper den ovanför en sökningscontainer.  
Om du samtidigt håller ned skifttangenten, så flyttas sökningen.  
Om det redan finns en sökning med samma namn, så öppnas dialogrutan Nytt namn där du först måste ange ett nytt namn för kopian som ska skapas.  
Om du drar sökningen till en sökningscontainer i stället för en tabellcontainer och släpper den där, så behandlas sökningen som en tabell.  
När du kopierar eller flyttar flera sökningar samtidigt genom att dra och släppa dem, kan du styra kopieringen för varje sökning separat.  
Nytt namn  
Här anger du ett nytt namn med vilket kopian ska sparas.  
När du vill flytta eller kopiera ett databasobjekt och det redan finns ett objekt med samma namn, så kan du ange ett namn med vilket kopian ska sparas i dialogrutan Nytt namn.  
Om du avbryter den här dialogrutan så startas kopieringen inte.  
Allmänt  
Här väljer du namn, typ och datakälla för databasen.  
I %PRODUCTNAME finns det flera olika sätt att arbeta med databaser:  
Du kan:  
integrera databaser i dBase - eller text -format i %PRODUCTNAME.  
komma åt en befintlig databas med ODBC eller JDBC.,  
komma åt en ADO -databas.  
Datakällan kan både vara en katalog i vilken det finns dBase-filer eller textfiler eller en datakälla i en befintlig databas som du vill ha åtkomst till.  
Vad du anger beror alltså på vilken datatyp som du vill registrera i %PRODUCTNAME.  
Adabas D-format  
Under Windows och Unix kan Adabas D-formatet användas.  
dBase - eller textformat  
Om du vill integrera filer i dBase - eller textformat behöver du inte göra så mycket mer än att ange den katalog där de här filerna finns.  
Varje fil listas då i databastabellen under fliken Tabeller så att de ska kunna integreras i %PRODUCTNAME som databastabeller.  
Åtkomst till externa databaser  
Även vid åtkomst till ett databassystem som erbjuder ett SQL-gränssnitt behöver du bara ange datakällan.  
I det här fallet rör det sig inte om en viss katalog, utan datakällan specificeras vanligen via sin beteckning.  
De är då så gott som direkt tillgängliga för dig när du arbetar i %PRODUCTNAME.  
Du får åtkomst till en extern SQL-databas via ODBC.  
Med ODBC kan du komma åt nästan vilken extern databas som helst som går att anropa med ODBC, under förutsättning att en passande ODBC-drivrutin är installerad.  
En ODBC-databas kan bara integreras om datorn har ett 32-bitars operativsystem och en 32-bitars ODBC-drivrutin.  
Namn  
Här anger du namnet med vilket du vill anropa databasen i %PRODUCTNAME.  
Det här namnet används bara för anrop av databasen i %PRODUCTNAME - det byts inte några namn på databasfiler.  
Förbindelse  
Databastyp  
Här anger du databastyp.  
Om du vill registrera en databas väljer du typ av databas bland databastyperna i kombinationsfältet.  
Du kan välja mellan typerna Adabas, dBase, Text, ODBC, JDBC, ADO, tabelldokument.  
URL för datakälla  
Här anger du den datakälla som du vill ha tillgång till som URL.  
Ett protokollschema placeras automatiskt framför, t.ex. "sdbc" eller "sdbc:dbase "elelr "jdbc".  
För databaser i Adabas-format anger du namnet på Adabas-filerna här.  
Om du har åtkomst till en extern Adabas-databas anger du datakällan så här: datornamn:databasnamn.  
Vid databaser i dBase - eller textformat utgör den katalog som innehåller dBase - eller textfilerna datakällan.  
I det här fallet anges här den kompletta sökvägen till respektive katalog.  
Men om du däremot vill få åtkomst till en extern databas, t.ex. via ODBC, anger du datakällan här.  
...  
Om du klickar på den här kommandoknappen öppnas en dialogruta där du kan välja en datakälla.  
För databaser av typen dBase eller Text kommer du till dialogrutan Välj ut sökväg där du väljer den katalog som innehåller din databas.  
Vid åtkomst till ODBC eller adressboksdrivrutinen öppnas dialogrutan Datakälla.  
Ny databas  
Den öppnar dialogrutan Skapa ny Adabas-databas.  
Datakälla  
Här väljer du den datakälla som du vill använda i %PRODUCTNAME.  
Om du vill registrera en extern databas i %PRODUCTNAME, måste du först ange datakällan i programmet.  
Datakällan omfattar både de data som användaren vill ha åtkomst till och den information som möjliggör åtkomsten till data.  
Om du vill ha åtkomst till en databas per ODBC, behöver du drivrutinen för den här databasen.  
Om den är installerad, så kan du definiera flera datakällor för varje installerad drivrutin.  
I den här dialogrutan visas de datakällor som är definierade för alla drivrutiner som finns installerade i systemet.  
Datakällor  
Här listas alla datakällor som du kan få åtkomst till.  
Förutom datakällans namn visas den tillhörande drivrutinen.  
Välj den datakälla som du vill registrera i %PRODUCTNAME.  
Administrera  
Med den här kommandoknappen öppnar du en dialogruta som kan vara olika för olika operativsystem och där du hanterar dina datakällor.  
Här kan du lägga till, radera eller konfigurera datakällor.  
Detta beskrivs i hjälpen till ditt operativsystem.  
ODBC  
Här gör du speciella inställningar för en databas som du får åtkomst till med ODBC.  
Till dessa räknas dina personliga åtkomstdata, eventuellt inställning av drivrutiner och definition av teckenuppsättning.  
En ODBC -databas finns för det mesta på en större dator i ett nätverk.  
Endast registrerade användare har åtkomst till den.  
En tabell måste ha ett entydigt index om du vill ändra eller lägga till dataposter i %PRODUCTNAME.  
ODBC-drivrutinerna är inte en del av %PRODUCTNAME. %PRODUCTNAME stöder bara ODBC 3 Standard.  
Användarnamn  
Här anger du ditt användarnamn för åtkomst till databasen.  
Lösenord krävs  
Markera den här rutan om det krävs ett lösenord för åtkomsten till databasen.  
Då efterfrågas alltid ditt lösenord när du ansluter till databasen första gången under en session.  
Drivrutinsinställningar  
I det här textfältet kan du, om du vill, ange ytterligare drivrutinsinställningar, i den mån det är nödvändigt.  
Teckenuppsättning  
Informationen som sådan ändras inte.  
DOS-baserade databaser använder i regel ASCII-teckenuppsättningen, som sammanfattas med olika kodsidor (landsspecifika teckenuppsättningar) under "IBMPC (850) / DOS ".  
Under Windows används teckenuppsättningen ANSI och Macintosh använder den teckenuppsättning som vi här kallar för "MAC".  
Om du anger "System" väljer du den teckenuppsättning som är standard för det operativsystem under vilket du har startat %PRODUCTNAME.  
Använd katalog för filbaserade databaser  
Om du markerar den här rutan används katalogen för den aktuella datakällan.  
Detta kan t.ex. vara nödvändigt om ODBC-datakällan är en databasserver.  
Men det kan uppstå problem vid användningen av katalog om ODBC-datakällan t.ex. är en dBase-drivrutin - i det här fallet bör du inte markera rutan.  
dBase  
Här gör du speciella inställningar för en dBase-databas.  
Med dBase menas här det speciella databas - och filformat som ursprungligen användes av Ashton Tates och senare Borlands databasprogram.  
Formatet betraktas som industristandard.  
Om det skrivs på annat sätt känns tabellerna inte igen.  
Visa inaktiva dataposter  
Markera alltid denna ruta när alla dataposter i filen ska visas, även sådana som markerats som raderade (inaktiva).  
Index  
I dialogrutan Index hanterar du indexen till dBase-tabellerna i den aktuella databasen.  
Index  
Här kan du hantera index till en dBase-databas.  
På det här sättet får du snabbare åtkomst till en databas om du söker data med hjälp av sorteringarna som är definierade genom index.  
När du skapar en tabell definierar du index på sidan med fliken Index.  
Tabell  
I den här listrutan väljer du önskad tabell.  
Tabellindex  
Om du vill ta bort ett eller alla index klickar du på kommandoknappen med motsvarande högerpil.  
Fria index  
I detta fält visas de fria index som för närvarande inte tilldelats någon tabell.  
Om du vill tilldela den valda tabellen ett index så markerar du det och klickar på vänsterpilen.  
Med den dubbla vänsterpilen tilldelar du tabellen alla fria index.  
<  
Om du klickar på den här ikonen överförs det markerade fria indexet till rutan Tabellindex.  
<<  
Om du klickar här överförs alla fria index till rutan Tabellindex.  
>  
Om du klickar på den här ikonen tas det markerade tabellindexet bort och överförs till rutan Fria index.  
>>  
Om du klickar på den här ikonen tas alla tabellindex bort och överförs till rutan Fria index.  
Text  
Här gör du speciella inställningar för import av en databas i textformat.  
Om en databas finns i textformat har informationen sparats som oformaterade ASCII-filer.  
I textformat finns varje post på en egen rad.  
Texterna i datafälten står för det mesta inom citattecken.  
Med textformat kan Du exportera innehållet från alla typer av databaser (även när det gäller ovanliga program och plattformar) och sedan importera denna information i ett annat program och på en annan plattform.  
Ett textexportfilter finns nästan alltid.  
Du kan använda %PRODUCTNAME Calc för att Redigera ASCII-filer eller databaser i textformat.  
Text innehåller sidhuvud  
Markera den här rutan om den första raden i filen innehåller fältnamnen.  
De tolkas då som kolumnhuvuden i databastabellen.  
Fältavgränsare  
Här anger du de tecken som används i filen för att skilja de enskilda datafälten åt.  
Du kan välja mellan följande tecken: semikolon (;), komma (,), kolon (:), tabb, blanksteg och ett eget tecken som du kan ange i kombinationsfältet.  
Textavgränsare  
Här anger du det tecken som identifierar textfält i databasen.  
Detta tecken får inte vara detsamma som fältavgränsaren.  
Om t.ex. citattecken ska användas som textavgränsare får det inte samtidigt vara fältavgränsare.  
Decimaltecken  
Här anger du den avgränsare som används för decimaltal.  
Beroende på de nationella inställningarna används komma (0,5) eller punkt (0.5).  
Tusentalsavgränsare  
Här anger du den avgränsare som används för tusental.  
Beroende på de nationella inställningarna används komma (1.000) eller punkt (1,000).  
Utökning  
I det här kombinationsfältet väljer du tillägget för textfilerna.  
Det valda tillägget bestämmer också delvis förinställningarna i de andra kombinationsfälten.  
Filnamnstillägget *.csv förutsätter att System anges som teckenuppsättning och att komma (;) anges som fältavgränsare.  
För filnamnstillägget *.sdf ändras dessutom teckenuppsättningen till "IBMPC (850) / DOS".  
Så här redigerar du en databastabell i textformat  
Men du kan importera tabellen till %PRODUCTNAME Calc, redigera den där och spara den med ett nytt namn som en databastabell i textformat.  
Öppna ett nytt tomt tabelldokument i %PRODUCTNAME Calc.  
Öppna datakällvyn, t.ex. genom att trycka på F4.  
Visa tabellen som du vill använda i datakällvyn.  
Klicka på kolumn - och radhuvudfältet uppe till vänster i datakällvyn för att markera hela tabellen.  
Släpp inte musknappen, utan dra tabellen direkt till det tomma tabellbladet i arbetsområdet.  
Släpp musknappen när du når fältet A1.  
Nu kan du redigera tabellens innehåll.  
Spara tabellen med kommandot Arkiv - Spara som och välj filtret "Text CSV" under Filtyp.  
Filemaker  
Här ställer du in Filemaker-databasens egenskaper.  
På en Macintosh kan du även importera det populära Filemaker-databasformatet till %PRODUCTNAME.  
Hämta alla dataposter på en gång  
Markera den här rutan om du vill importera samtliga dataposter i Filemaker-filen.  
Maximalt antal dataposter  
Om du har aktiverat Hämta alla dataposter på en gång kan du begränsa antalet dataposter som ska hämtas samtidigt här (gäller mycket stora databaser).  
Administrera datakällor  
Här öppnas en dialogruta där du kan administrera datakällor i %PRODUCTNAME.  
Till vänster i dialogrutan finns det en lista över registrerade datakällor.  
Varje datakälla i listan visar sin status med en symbol:  
oförandrad  
markerad för radering  
markerad som ny databas  
markerad för ändring av egenskaper  
Om du avslutar dialogrutan med OK eller klickar på Använd utförs de markerade ändringarna.  
Om du avslutar dialogrutan med Avbryt görs inga ändringar.  
Varje namn på en datakälla får bara förekomma en gång.  
Det enda undantaget från den här regeln gäller en datakälla som har markerats för radering: du får använda den datakällans namn till en ny datakälla.  
Du registrerar en ny datakälla genom att klicka på kommandoknappen Ny datakälla eller med kommandot Ny datakälla på snabbmenyn.  
Du kan radera posten i listan på postens snabbmeny:  
Radera datakälla.  
Med hjälp av kommandot Återställ datakälla på snabbmenyn till en datakälla som är markerad för radering kan du ångra detta.  
I dialogrutan finns följande flikar som alltid relaterar till den databas som är markerad i listan till vänster:  
Under fliken Allmänt kan du välja en Databastyp.  
Beroende på vad du väljer finns det sedan en ytterligare flik med Namnet på databastypen (se följande hyperlänkar).  
Posten Tabelldokument är ett undantag; det finns ingen egen flik för den.  
Dessutom finns flikarna Tabeller, Sökningar och Länkar.  
Beroende på vilken typ av databas som du väljer visas någon av följande flikar:  
Tabelldokument  
Med den här databastypen väljer du ett tabelldokument från %PRODUCTNAME Calc eller MS Excel som datakälla.  
Under fliken Tabeller kan du välja bland alla tabeller som inte är tomma och inte är dolda i dokumentet.  
Om du vill använda en hel tabell som datakälla måste data börja i cell A1; på rad 1 måste det stå kolumnrubriker.  
Om dataområden har definierats i tabelldokumentet kan du välja varje dataområde som egen databastabell.  
Det går bara att läsa data, inte att skriva data.  
Utföra SQL-sats  
Med kommandot SQL på snabbmenyn till en databas öppnas en dialogruta där du kan mata in ett SQL-kommando för administration av databasen direkt.  
Kommandot leder inte till att något filtrerat databasinnehåll visas; dialogrutan är bara till för att mata in administrationskommandon som t.ex. Grant (tilldela användarbehörighet), Create Table (skapa tabell), Drop Table (radera tabell) och så vidare.  
Datakällan måste stödja SQL-kommandona - dBase kan t.ex. inte utföra alla kommandon som nämns här.  
I ett särskilt statusfönster visas om kommandot verkställs som det ska.  
Om du vill utföra en SQL-sökning för att filtrera data från en databas, öppnar du Sökningsutkast.  
Kommando att utföra  
Här skriver du SQL-instruktionen.  
I den öppnade datakällan "Bibliography" kan du t.ex. ange följande SQL-kommando:  
SELECT "Address" FROM "biblio ""biblio"  
Om du vill ha utförligare information om SQL-kommandon bör du läsa litteratur i detta ämne.  
Föregående kommandon  
Här visas de föregående kommandona.  
Om du markerar ett kommando överförs det till fältet Kommando att utföra.  
Status  
Här visas statusuppgifter för SQL-databasen som visas efter att SQL-kommandot har utförts.  
Om det finns fel i SQL-syntaxen får du information om var felet finns.  
Utför  
Klicka på Utför när du vill starta kommandot.  
Tabeller  
Här är alla tabeller som hör till den aktuella databasen listade.  
I listrutan väljer du vilka tabeller som ska visas i %PRODUCTNAME genom att klicka med musen på de tillhörande kryssrutorna.  
Dessutom går det att redigera tabellstrukturen, definiera nya tabeller och radera tabeller.  
Tabeller från databaser som stöder "Catalog" eller "Schema "visas i en hierarkisk vy.  
Du kan sortera tabeller med hjälp av snabbmenyn.  
Nytt tabellutkast  
Öppnar Tabellutkast -fönstret där du kan skapa en ny tabell.  
Redigera tabell  
Öppnar Tabellutkast -fönstret där du kan redigera den markerade tabellen.  
Radera tabell  
Raderar den markerade tabellen efter en säkerhetskontroll.  
Filter  
Här bestämmer du vilka tabeller som ska visas i %PRODUCTNAME.  
Du markerar tabellerna i listrutan Filter.  
Om du markerar en överordnad post visas posten i fetstil och alla underordnade poster markeras automatiskt.  
Detta gäller också om t.ex. en tabell tillkommer genom att en fil kopieras: även den markeras.  
Om du bara markerar alla underordnade poster som är synliga visas den överordnade posten inte i fetstil.  
Det betyder t.ex. att tabeller som läggs till i efterhand inte är markerade till att börja med.  
Visa versionskolumner (om tillgängliga)  
En del databaser, t.ex. Adabas, har ett internt datafält med ett versionsnummer för varje datapost.  
Om dataposten ändras höjs versionsnumret med 1.  
Om du har markerat den här rutan kan du se det interna versionsnumret på dataposten i databastabellen.  
På snabbmenyn till tabeller finns följande kommandon:  
Sortera stigande  
Sorterar tabellen efter namn i stigande alfabetisk ordning.  
Sortera fallande  
Sorterar tabellen efter namn i fallande alfabetisk ordning.  
JDBC  
Här gör du speciella inställningar för en databas som du har åtkomst till via JDBC.  
Drivrutinsklasserna måste anges i filen java.ini eller under Verktyg - Alternativ - %PRODUCTNAME - Säkerhet i fältet ClassPath.  
JDBC-drivrutinsklass  
För uppkopplingen mot databasen behövs en JDBC-drivrutin som du måste ange här.  
URL  
Ange t.ex. "jdbc:mysql: / /<servernamn> / <DB-namn>" för en MySql-JDBC-drivrutin, där "servernamn "är serverns namn och DB-namn är databasen namn.  
För en närmare beskrivning för din drivrutin hänvisar vi till dokumentationen för drivrutinen.  
Adabas D  
Här loggar du in dig för en databas i Adabas-format.  
För att kunna göra detta måste du ange användarnamn och lösenord.  
Mer information om databasformatet Adabas D.  
Användarnamnet får bestå av högst 18 tecken.  
Lösenordet måste vara minst 3 och högst 18 tecken långt.  
Användarinställningar  
Här administrerar du användarna av en Adabas - eller ADO-databas.  
Mer information om databasformatet Adabas D.  
Användarurval  
Användare  
Här markerar du användaren vars inställningar du vill administrera.  
Lägg till användare  
Klicka här om du vill lägga till en ny användare för den här datakällan.  
Ändra lösenord  
Här ändrar du lösenordet för en markerad användare för den här datakällan.  
Radera användare  
Här raderar du en markerad användare.  
Åtkomsträttigheter för markerad användare  
Här ser och redigerar du åtkomsträttigheterna för en markerad användare.  
Om fälten inte är aktiverade har du inte rättighet att ändra rättigheter för den markerade användaren.  
ADO  
Här registrerar du en databas i formatet ADO (Microsoft ActiveX Data Objects), bl.a. för åtkomst till MS Access-databaser.  
Du anger URL och användarnamn och definierar om ett lösenord behövs.  
För att du ska kunna använda ADO måste Access 2000 eller uppdateringen från www.microsoft.com / data vara installerad.  
URL  
Här anger du URL.  
PROVIDER=Microsoft.Jet.OLEDB.4.0; DATA SOURCE=c:\Access\nwind2000.mdb  
Det här exemplet visar en koppling till en Access 2000-fil.  
DSN=SQLSERVER  
Det här exemplet använder ODBC-drivrutinen som provider.  
Användarnamnet får bestå av högst 18 tecken.  
Lösenordet måste vara minst 3 och högst 18 tecken långt.  
Statistik Adabas D  
Här definieras åtkomstalternativ för administrationen av en lokal databas i Adabas-format.  
Här kan administratören tilldela särskilda behörigheter för ändringar av tabeller i respektive tabells dialogruta för egenskaper.  
Databuffertstorlek  
Här kan du ändra storleken på databasens databuffert (den virtuella minnesförbrukningen).  
Den nya storleken är tillgänglig när databasen har startats om.  
Tillväxtstorlek  
Här ändrar du tillväxtstorleken, som är den storlek med vilken databasen automatiskt utökas när den är för liten för att ta emot nya data.  
Den nya storleken är tillgänglig när databasen har startats om.  
Den databas som följer med %PRODUCTNAME är begränsad till 100 MB.  
Användarnamn Control  
Här anger du namnet på Control-användaren.  
Lösenord Control  
Här anger du Control-användarens lösenord.  
Stäng service när %PRODUCTNAME avslutas  
Om den här rutan är markerad, avslutas Adabas-databasservern när du avslutar %PRODUCTNAME.  
Detta gäller bara om databasservern har startats från %PRODUCTNAME och om Control-användaren har angetts med lösenord.  
Utvidgat  
Här öppnar du dialogrutan Databasstatistiker.  
Databasstatistiker  
För en databas i Adabas-format visas här statistiska uppgifter; bland annat hur många procent av databasens minnesutrymme som används.  
Databasfiler  
SYSDEVSPACE  
Här visas sökväg och namn för SYSDEVSPACE.  
TRANSACTIONLOG  
Här visas sökväg och namn för filen TRANSACTIONLOG.  
DATADEVSPACE  
Här visas sökväg och namn för filen DATADEVSPACE.  
Databasstorlekar  
Totalstorlek (MB)  
Här anges den totala storleken (i megabyte).  
Fritt minne (MB)  
Här anges det lediga minnesutrymmet (i megabyte).  
Minnesutnyttjande (i%)  
Här anges hur många procent av den totala storlekens minnesutrymme som är upptaget.  
Sökningar  
Här listas alla sökningar som hör till den aktuella databasen.  
Du kan bara öppna den här fliken för en ny datakälla om du har sparat ändringarna i dialogrutan Verktyg - Datakällor innan.  
En dialogruta informerar dig eventuellt om detta och ger dig möjlighet att spara.  
Sökningar  
I listrutan administrerar och startar du sökningarna för den aktuella datakällan.  
Nytt sökningsutkast  
Här skapar du en ny sökning.  
Fönstret Sökningsutkast visas.  
Mata in nytt SQL-kommando  
Öppnar ett fönster där du kan mata in en ny sökning per SQL.  
Redigera sökning  
Här redigerar du en markerad sökning.  
Fönstret Sökningsutkast visas.  
Mata in SQL-kommando  
Öppnar ett fönster där du kan redigera den aktuella sökningen på SQL-språk.  
Radera sökning  
Här raderar du en markerad sökning.  
Byt namn  
Öppnar dialogrutan Klistra in som.  
Namn på sökning  
Ange sökningens namn.  
Länkar  
Här listas alla angivna länkar till formulärdokument för den aktuella datakällan.  
Formulär och länkar  
I %PRODUCTNAME har du tillgång till datakällorna som du registrerar och administrerar under Verktyg - Datakällor.  
I datakällvyn (F4) visas data i tabellform till höger och till vänster, i Explorer för datakällor, datakällorna med deras länkar, sökningar och tabeller.  
Du kan tilldela dina dokument, t.ex. textdokument eller tabelldokument, en datakälla som Länk.  
Detta används bara för att få en snabb tillgång till dokument från datakällvyn - en ytterligare länk mellan dokument och datakälla är visserligen möjlig, men inte nödvändig.  
I dina dokument, oberoende av om du skapar en länk eller inte, kan du också använda fältkommandon fältkommandon och / eller formulärfunktioner och referera till respektive aktuellt innehåll i en datakällas datafält.  
Med formulärfunktionerna kan du till exempel skapa formulär.  
Alla text - eller tabelldokumenten kan ha innehåll från datakällor.  
De här och andra dokument kan du lägga till som länk i datakällvyn, för att lättare få tillgång till de här dokumenten från datakällvyn.  
Du måste själv administrera de här länkarna.  
Länkar  
I listrutan administrerar du länkarna för den aktuella datakällan.  
Ny länk  
Här skapara du en ny länk.  
Dialogrutan Dokumentlänk - ny visas:  
Namn  
Ange namnet på länken här.  
URL  
Ange URL:en eller klicka på... och välj den.  
Redigera länk  
Här redigerar du en markerad länk.  
Dialogrutan Dokumentlänk - redigera visas som motsvarar dialogrutan Dokumentlänk - ny.  
Radera länk  
Här raderar du en markerad länk.  
Det är bara tilldelningen av det här dokumentet till datakällan som raderas, inte själva dokumentet.  
Öppna dokument  
Dokumentet är skrivskyddat när det öppnas.  
Redigera dokument  
Öppnar det angivna dokumentet i en markerad länk för redigering.  
Nytt formulär  
Öppnar ett nytt dokument av den valda dokumenttypen.  
Foga in formulärfält eller fältkommandon om du vill och spara dokumentet.  
Det förs automatiskt in som länk.  
LDAP  
Här gör du inställningar för en LDAP-server som du har registrerat som databastyp Adressbok.  
Värddatornamn  
Här anger du namnet på LDAP-servern, t.ex.: ldap.server.com.  
Base DN  
Här anger du ytterligare parametrar som LDAP-servern behöver, t.ex.: dc=com.  
Portnummer  
Här anger du LDAP-serverns portnummer, t.ex. 389.  
Dataposter (max)  
Här anger du hur många dataposter som maximalt laddas vid åtkomst till LDAP-servern.  
Adabas D-databas  
Med %PRODUCTNAME levereras en något förminskad version.  
Närmare information om Adabas, fler hjälpfiler samt möjlighet att beställa senare versioner finns hos tillverkaren på adressen http: / /www.adabas.com.  
Du måste kunna nå Adabas-databasservern för att kunna arbeta med en Adabas-databas.  
Om du inte använder en Adabas-databasserver i nätverket utan t.ex. arbetar på en fristående dator, måste du först installera och starta serverprogrammet.  
Det serverprogram som medföljer %PRODUCTNAME kan installeras med ett särskilt setupprogram.  
Setupprogrammet för installation av Adabas D startar automatiskt efter setupprogrammet för %PRODUCTNAME om du gör en fristående installation.  
Det finns mer information om Adabas-installationen i det separata installationsdokumentet.  
Egenskaper hos %PRODUCTNAME -versionen av Adabas  
Adabas D, version 11, som medföljer %PRODUCTNAME, är begränsad till databasstorleken 100 MB.  
Vid användning i nätverk kan högst tre användare samtidigt komma åt databasen.  
Det finns mer information i filen license.txt som finns i Adabas-katalogen efter installationen.  
Adabas bör inte installeras i %PRODUCTNAME -katalogen utan i en egen katalog.  
Adabas och %PRODUCTNAME kan avinstalleras oberoende av varandra.  
Vid installationen aktiveras bl.a. miljövariabeln DBROOT, som hänvisar till den katalog där du har installerat Adabas.  
Det innebär att du måste starta om datorn innan du använder Adabas för första gången.  
Om miljövariabeln DBROOT hittas vid installationen kan du inte installera Adabas, eftersom setupprogrammet i så fall utgår ifrån att en Adabas-version redan har installerats.  
Du kan också använda SQL-kommandon för att administrera den.  
I %PRODUCTNAME stöder Adabas kommandon enligt standarden SQL92.  
Prestanda för Adabas D i %PRODUCTNAME  
%PRODUCTNAME kan ha åtkomst till en Adabas D-databas, om det är version 11.02 eller högre.  
För Adabas D-versionen 11 i %PRODUCTNAME gäller följande värden:  
Begränsning till 100 MB och 3 användare per databas.  
Adabas D stöder följande datatyper:  
Datatyp  
Innehåll  
CHAR (N) N <= 254  
Teckensträngar i ASCII - eller EBCDIC-kod eller som BYTE.  
VARCHAR (N) N <= 254  
Den interna arkiveringen av CHAR-värden görs upp till en längd av 30 tecken i fast format.  
Större CHAR-värden lagras alltid internt med variabel längd.  
Genom användning av datatypen VARCHAR kan även CHAR-värden med en längd under 30 lagras med variabel längd.  
BOOLEAN  
För att skilja mellan "finns / finns inte" och "sant / falskt ".  
DATE  
Lagras som internt format YYYYMMDD.  
Den externa visningen kan konfigureras.  
TIME  
TIME-värden lagras internt på formen HHMMSS.  
Liksom med DATE-värden går det att konfigurera den externa visningen.  
DATE - och TIME-värden är speciella CHAR-värden.  
Det betyder att utöver datum - och klockslagsfunktionerna kan även alla funktioner för CHAR-värden användas.  
TIMESTAMP  
TIMESTAMP-värden lagras internt på formen ÅÅÅÅMMDDTTMMSSmmmuuu.  
De utgör en kombination av ett DATE - och ett TIME-värde och är utvidgade till att ange milli - och mikrosekunder.  
Förutom användningen som tidsstämpel kan TIMESTAMP-värden även användas för tidsberäkning, eftersom övergång till nästa dag därvid inte behöver behandlas av användaren.  
TIMESTAMP-värden är speciella CHAR-värden.  
Det betyder att utöver datum - och klockslagsfunktionerna kan även alla funktioner för CHAR-värden användas.  
FIXED (N,M)  
För numeriska värden innebär detta en lagring med högst 18 positioner och fast decimalkommaplacering.  
FLOAT (N)  
En decimal flyttalslagring med maximal noggrannhet på 18 positioner.  
LONG  
För lagring av oformaterade data (BLOBs) finns i Adabas datatypen LONG, som kan ta emot upp till 2,1 GB data per kolumn.  
Liksom för CHAR-kolumner stöds varianterna ASCII, EBCDIC och BYTE.  
Därmed kan Adabas organisera omfångsrika text-, bild - och ljuddata på lämpligt sätt.  
De ytterligare datatyper som förekommer i SQLMODE tolkas av Adabas och avbildas på ovan angivna datatyper.  
Skapa ny Adabas-databas  
I dialogrutan Skapa ny Adabas-databas kan du skapa en ny Adabas-databas.  
Den här dialogrutan kan du t.ex. öppna på följande sätt:  
Öppna dialogrutan Administrera datakällor via Verktyg - Datakällor.  
I fältet Databastyp väljer du datatypen "Adabas".  
Klicka på kommandoknappen Ny databas.  
I %PRODUCTNAME är flera fält i dialogrutan redan ifyllda, och du behöver normalt bara ange databasens namn samt administratörens namn och lösenord.  
De här tre uppgifterna är obligatoriska.  
Radera Adabas-databas  
Om du raderar databasposten i %PRODUCTNAME, raderar du enbart åtkomsten till informationen från %PRODUCTNAME.  
De "egentliga" filerna i databasen finns kvar.  
Om du verkligen vill radera alla filer, gör du så här:  
Ange databasens namn. (Det är inte nödvändigtvis samma namn som visas på posten.) Välj Egenskaper.  
Under fliken Typ står databasens namn i fältet Datakälla.  
Ta reda på vilka mappar systemvariablerna DBCONFIG och DBWORK pekar på.  
I Unix definieras de här variablerna i ett Startscript.  
I katalogen $DBCONFIG$ raderar du tre filer med databasens namn.  
Om din databas t.ex. heter TEST, raderar du följande filer vid en typisk installation under Windows:  
C:\Adabas\Sql\Test.sys, Test.trs och Test.dat.  
I katalogen $DBCONFIG$\Config raderar du en fil med databasens namn.  
Om din databas t.ex. heter TEST raderar du filen C:\Adabas\Sql\Config\Test.  
I katalogen $DBWORK$\Wrk raderar du en komplett katalog med databasens namn.  
Om din databas t.ex. heter TEST raderar du katalogen C:\Adabas\Sql\Wrk\Test.  
Var noga med att bara radera de filer och den mapp som har samma namn som databasen.  
Manuell start och avstängning av en Adabas-databas  
NoDBService  
ställer databasen på COLD.  
xutil -d <DBNAME> -u <CONTROLUSER>,<CONTROLPASSWORT> shutdown  
ställer databasen på COLD.  
xutil -d <DBNAME> -u <CONTROLUSER>,<CONTROLPASSWORT> restart  
ställer databasen på WARM.  
stp -d <DBNAME> -NoDBService  
stänger av databasen helt och hållet.  
Felmeddelanden för en Adabas-databas  
Nedan beskrivs några felmeddelanden som kan uppträda vid arbetet med Adabas D.  
Databasen kan inte stängas av / startas om så länge någon användare är ansluten till den.  
Stänga alla aktiviteter som eventuellt fortfarande är öppna och som visar det här databasinnehållet.  
Vid fleranvändarsystem måste du be alla användare att lämna databasen.  
Om detta inte hjälper måste du även avsluta %PRODUCTNAME och sedan starta om.  
Client unable to establish connection; -813 SERVERDB MUST BE RESTARTED  
Det här felet uppstår om du försöker komma in i en Adabas D-databas som inte har startats.  
Men då måste Control-användaren vara definierad i databasens egenskaper.  
Detta görs när databasen skapas.  
Client unable to establish connection; -8022 USER ALREADY CONNECTED  
Det här felet uppstår om du försöker komma in i en Adabas D-databas, men samma användare redan är ansluten till databasen.  
Fel vid skrivning av data i databasen  
"Databasens egenskaper kan inte ändras eftersom databasen fortfarande används." Om du ser det här felmeddelandet måste du avsluta och starta om %PRODUCTNAME.  
Sedan ändrar du direkt databasens egenskaper.  
Adabas-server i nätverk  
Om användningen av databasen är delad i ett nätverk, körs Adabas-servern i nätverksdatorn medan enbart klienten körs i arbetsstationerna.  
Remote Connection  
För att en "Remote connection" (fjärranslutning) ska vara möjlig, måste hjälpprogrammet xtcpupd.exe köras på båda datorerna (klient och server).  
Programmet xtcpupd.exe finns bara för Windows.  
På servern måste programmet x_server från katalogen adabas / bin Adabas / bin startas (alla plattformar).  
Du registrerar en fjärranslutning (remote connection) som ny Adabas-databas.  
I textfältet Datakälla matar du in namnet på den externa datorn, ett kolon och namnet på den externa databasen, t.ex. datornamn:databas.  
Ange användarnamn och lösenord under fliken Adabas D och klicka på OK.  
Nu kan du använda fjärrdatabasen.  
Om du vill skapa en ny databas på en fjärrserver, finns det två möjligheter:  
Du kan installera %PRODUCTNAME på fjärrservern och skapa den nya databasen (lokalt) där, eller  
Du kan använda Adabas-verktygen till att skapa en ny Adabas-databas på servern.  
Det är inte möjligt att skapa den nya databasen från en %PRODUCTNAME -klient.  
Skapa ny Adabas-databas  
I den här dialogrutan skapar du en ny Adabas-databas.  
Databasnamn  
Här anger du namnet på databasen i Adabas.  
Användarinställningar  
Här gör du användarinställningarna. %PRODUCTNAME har fyllt i fälten så långt som möjligt med lämpliga förinställningar.  
Administratör  
Här anger du namnet på databasens administratör.  
När en ny Adabas-databas skapas, måste du ange minst ett administratörsnamn och ett tillhörande lösenord.  
Administratören är även den första användaren.  
Den Adabas-version som medföljer %PRODUCTNAME tillåter tre samtidiga användare.  
Det här fältet visas bara om du öppnar dialogrutan via Ny datakälla.  
Control-användare  
Control-användaren har behörighet att ändra parametrar i databasen.  
Normalt lämnar du control-användarens förinställda namn och lösenord oförändrade.  
Control-användaren berörs inte av begränsningen till tre användare.  
Domän-användare  
En domänanvändare måste finnas internt i Adabas.  
Normalt lämnar du domänanvändarens förinställda namn och lösenord oförändrade.  
Domänanvändaren berörs inte av begränsningen till tre användare.  
Det här fältet visas bara om du öppnar dialogrutan via Ny datakälla....  
Lösenord  
Det används även automatiskt för både control-användaren och domänanvändaren.  
Du kan även använda olika lösenord om du vill.  
Databasinställningar  
Här gör du databasinställningarna. %PRODUCTNAME har fyllt i fälten så långt möjligt med lämpliga förinställningar.  
DEVSPACEs är enheter eller filer som innehåller delar av Serverdb.  
För Adabas rekommenderar vi att du lagrar var och en av de olika DEVSPACE på var sin hårddisk.  
Sökvägarna till filerna inklusive filnamn får inte bestå av mer än 40 tecken.  
SYSDEVSPACE  
Ange adressen till System Devspace här.  
I denna Devspace lagras bl a konfigurationsdata.  
Dess storlek är direkt proportionell mot databasens storlek.  
TRANSACTIONLOG  
Ange här adressen till transaktionsloggfilen.  
Ändringar i datauppsättningen registreras i loggen och kopieras vid transaktionens slut.  
Transaktionsloggen är till för att möjliggöra rollback (återföring av transaktioner) och fylls i cykliskt.  
Den måste vara tillräckligt stor för att rymma ändringar av alla öppna transaktioner.  
DATADEVSPACE  
Ange här adressen till Data Devspaces.  
Där lagras användardata (tabeller, index) och SQL-katalogen (Schema Information).  
De data som hör till en tabell fördelas likformigt av Adabas på alla Data Devspaces.  
Det diskutrymme som definieras av alla Data Devspaces utgör databasens fulla storlek.  
I %PRODUCTNAME -versionen av Adabas är det utrymmet begränsat till 100 MB per databas.  
Om du behöver större kapacitet bör du vända dig till Adabas tillverkare, Software AG, på adressen www.adabas.com.  
Om alla Data Devspaces är fyllda till 100%, avbryts driften av databasen och en "Emergency Shutdown" (nödstopp) inträffar.  
Databasen förstoras därpå automatiskt med ett inkrementvärde (upp till 100 MB) och startas om.  
Denna åtgärd innebär att sparad information inte förstörs.  
...  
Här öppnar du en dialogruta där du kan spara Adabas-systemfilen för den aktuella databasen.  
Välj en katalog och ange namnet.  
Transaktionsfil (MB)  
Här väljer du storlek (i MB) för transaktionsfilen.  
Databasstorlek (MB)  
Här väljer du storlek (i MB) för databasen.  
I %PRODUCTNAME -versionen är den begränsad till 100 MB.  
Databuffertstorlek (MB)  
Här väljer du storlek (i MB) för databufferten (datacachen).  
I den här cachen finns de sidor i Data Devspaces där den senaste läsningen eller skrivningen gjordes.  
Den används gemensamt av alla samtidiga användare.  
Träffkvoten, d.v.s. förhållandet mellan lyckade och misslyckade sökningar i cachen, är av avgörande betydelse för prestandan. (Med en lyckad sökning menas att den sökta informationen hittas i cachen.)  
Allmänt  
Under den här fliken listas allmänna egenskaper för det aktuella objektet.  
Till dessa egenskaper hör både det namn som du kan ange eller ändra för vissa objekt och diverse information om objektet.  
Därför visas bara den information och det innehåll som är relevant för objektet ifråga.  
Namn  
I textfältet anges det namn med vilket objektet visas.  
Om objektet ännu inte fått något namn skriver du ett här.  
För en del objekt kan du även ändra de namn som objekten tilldelats.  
När du registrerar en databas anger du här det namn under vilket den ska registreras i %PRODUCTNAME.  
Du kan ange vilket namn du vill, men vissa tecken är inte tillåtna (t.ex. /,\,?, #) och ignoreras när du försöker skriva dem.  
När du väljer namn gäller bara filsystetmets begränsningar som är specifika för operativsystemet.  
Om Du arbetar i ett nätverk bör Du tänka på att namnen på de lokala databaserna inte får vara identiska med namn på databaser på en nätverksserver.  
Om Du t ex vill lägga upp ett nytt formulär för en databas på en nätverksserver kan %PRODUCTNAME bara skapa en referens till denna databas om det inte finns en databas med samma namn på Din lokala hårddisk.  
Skrivskyddad  
Markera den här rutan om du vill skrivskydda filen.  
Den är då bättre skyddad mot oavsiktliga ändringar och raderingar.  
Avmarkera rutan om du vill kunna skriva över eller radera en fil.  
Den här kryssrutan visas när du tittar på en fils egenskaper, det vill säga när du t.ex. undersöker den i en mapp.  
Den här rutan visas inte i egenskapsdialogrutan i ett öppnat dokument.  
Ytterligare information  
Denna ytterligare information kan Du visa, dölja, inskränka till vissa dokumentegenskaper eller utöka med mer information.  
Här presenteras all information, oberoende av om en mapp, en databas eller något annat har markerats:  
Typ  
Det kan t.ex. röra sig om en fil, en länk eller en speciell databastyp.  
Beroende på typ anges dessutom följande data:  
Plats  
Här ser Du den kompletta sökvägen till objektet.  
Storlek  
Här anges objektets storlek i byte, kB eller MB.  
Antal innehåll  
Om Gallery är markerat visas antalet teman.  
Skapat  
Även namnet på den som skapat objektet anges.  
Ändrat  
Här anges även namnet på den som gjort ändringen.  
Utskrivet:  
Här anges datum och klockslag för den senaste utskriften.  
Version:  
Här anges dokumentets versionsnummer.  
Mall:  
Om Du har använt en dokumentmall anges namnet på mallen här.  
Redigeringstid:  
Den totala redigeringtiden fram tills nu anges här.  
Här väljer du symbolvy av Gallery-temat.  
Här väljer du detaljvy av Gallery-temat.  
Gallery  
Här öppnar du Gallery, grafik - och ljudhanteringen i %PRODUCTNAME.  
Du kan lägga till fler grafikobjekt, ljud och teman.  
Till vänster ser du teman.  
För varje tema som du klickar på, visas objekten som det innehåller till höger.  
Du kopierar bilder mellan Gallery och dokument med dra-och-släpp.  
Objekten kan visas som symboler (symbolvy) eller i en lista (detaljvy).  
Om du dubbelklickar på ett objekt eller på blanksteg byter du mellan visning av flera objekt och ett enda objekt.  
Så här lägger du till ett nytt tema till Gallery.  
Klicka på kommandoknappen Nytt tema.  
Nu öppnas dialogrutan Egenskaper för Nytt tema med flikarna Allmänt och Filer.  
Om du har lagt till en extra Gallery-sökväg under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar, kan du bara redigera Gallery-teman via denna extra sökväg.  
Via den extra sökvägen kan du däremot skapa, redigera och radera dina egna teman.  
Nytt tema  
Med den här kommandoknappen lägger du till ett nytt tema till Gallery.  
Dialogrutan Egenskaper för Nytt tema visas.  
Ange ett namn för temat under fliken Allmänt och lägg till nya filer under fliken Filer.  
Du kan också välja Egenskaper på temats snabbmeny till vänster i Gallery -fönstret och lägga till nya filer under fliken Filer.  
Du kan välja bland följande poster på snabbmenyerna:  
Egenskaper  
Det här kommandot öppnar dialogrutan Egenskaper för (tema) för ett markerat tema i Gallery.  
Det finns följande flikar:  
Filer  
Ljudservrar som stöds  
Om du vill kunna använda ljudfunktionerna, så måste programvaran Network Audio System från NCD Inc. vara installerad på den dator på vilken ljudet ska spelas (och givetvis krävs ljud-hårdvara som stöds).  
Det finns även att hämta på andra webbsidor.  
Du behöver version 1.2 pl 4 eller högre.  
Men vissa tillverkare bifogar inte NAS!  
För närvarande stöds följande system av NAS:  
Linux x86 (om det finns ljuddrivrutiner för kortet - sådana finns dock för nästan alla kort), SGI, HP, SUN.  
Detta gäller bara för ljudservern, d.v.s. den dator som ska låta spela upp ljuden, "den med högtalarna".  
Klienterna (d.v.s. %PRODUCTNAME -programmen) berörs inte alls av detta, de kan kommunicera med vilken NAS-ljudserver som helst, oavsett på vilken hårdvara den körs.  
Formatet är likadant som för DISPLAY-variabeln, t ex name:0  
Ifall AUDIOSERVER inte har angetts, så används DISPLAY-variabeln (sedan är alltså ljud och video på samma dator).  
Ifall DISPLAY-variabeln inte heller har angetts (därför att bildskärmen t ex har angetts via kommandoraden), så fungerar inte ljudet. (Ljudservern kan alltså inte anges via kommandoraden.)  
Du kan även använda rplayd för att spela upp ljud.  
Men bara en ljudserver kan vara aktiv.  
När du arbetar med rplayd kan du t.ex. inte längre lyssna på ljud under KDE eftersom KDE använder sin egen ljudserver.  
Du bör helst starta rplayd innan X Window startas.  
Dessutom kan du med SalSound och OSS (Open Sound System) spela upp ljud på den lokala displayen.  
Så småningom ska det även gå att spela upp *.au - och *.snd-filer.  
Filer  
Här lägger du till nya filer till det markerade temat.  
Filtyp  
Välj den filtyp som ska sökas.  
Hittade filer  
I denna flerradiga listruta visas sökresultatet.  
Du kan markera enstaka påträffade filer och lägga till dem till det aktuella temat med kommandoknappen Lägg till.  
Dessutom kan Du använda tangenterna Skift och Kommando Ctrl för att välja ut sammanhängande eller uppdelade områden med filer i listan.  
Sök filer...  
Klicka på den här knappen om Du vill öppna en urvalsdialog för mappar.  
Här väljer Du den mapp, där Du vill söka.  
Dialogrutan innehåller även kryssrutan Undermappar.  
Undermappar  
Markera detta fält i mapp-urvalsdialogen om Du även vill att den valda mappens alla undermappar ska genomsökas.  
Lägg till  
Om Du klickar på den här knappen adderas alla markerade filer till det valda temat.  
Filerna kopieras inte, utan infogas endast som referenser i Gallery.  
Lägg till alla  
Om Du klickar på den här knappen adderas alla påträffade filer till det valda temat.  
Filerna kopieras inte, utan infogas endast som referenser i Gallery.  
Förhandsvisning  
Markera detta fält om Du vill se en förhandsvisning av varje hittad fil när Du klickar på den.  
Förhandsvisningsfält  
Här ser du en förhandsvisning av den markerade filen.  
Första steg  
Så här kan du underlätta arbetet med hjälp av våra exempel - och dokumentmallar.  
Med %PRODUCTNAME får du ett stort antal exempeldokument och dokumentmallar.  
Du öppnar dem via Arkiv - Nytt - Mallar och dokument eller via tangentkombinationen Skift + Kommando Ctrl +N.  
När du öppnar en av dokumentmallarna, skapas ett nytt namnlöst dokument som baserar på den här mallen.  
Ett flertal AutoPiloter (i meny Arkiv) hjälper dig att skapa egna skräddarsydda dokumentmallar, t.ex. för brev, fax, presentationer eller webbsidor som du sedan kan använda som grund för dina andra dokument.  
Använd de medföljande dokumentmallarna direkt eller för att lära dig tekniker när du arbetar med %PRODUCTNAME.  
Om du utformar en tidning, skriver en bok, ordnar din ekonomi, eller vill göra formulär och avtal eller ett cd-omslag, är chansen ganska stor att %PRODUCTNAME redan innehåller dokumentmallar för de här och många andra uppgifter!  
Arbeta med %PRODUCTNAME  
Arbeta med textdokument  
Arbeta med tabelldokument  
Arbeta med presentationer  
Arbeta med teckningar  
Arbeta med formler  
Sätta på / stänga av aktiv hjälp  
Den aktiva hjälpen visar förutom funktionsnamnet en kort funktionsbeskrivning när du placerar markören på en kommandoknapp, ett annat kontrollfält eller en ikon.  
Så sätter du på och stänger av den aktiva hjälpen:  
Klicka på Hjälp på menyraden i programmet och välj Aktiv hjälp.  
En bock bredvid menyposten visar att den aktiva hjälpen är aktiverad.  
Så här aktiverar du den aktiva hjälpen temporärt:  
Tryck på tangentkombinationen Skift+F1 för att aktivera den aktiva hjälpen.  
Muspekaren visar ett frågetecken.  
Du kan föra den här Hjälpmuspekaren över alla kontrollelement, ikoner och menypunkter och få lite information om respektive kommando.  
Nästa gång du klickar med musen inaktiveras Hjälpmuspekaren igen.  
Inaktivera URL-igenkänning med AutoKorrigering  
När du skriver text känner %PRODUCTNAME automatiskt igen om ordet kan vara en URL och ersätter det här ordet med en hyperlänk. %PRODUCTNAME formaterar hyperlänken med direkta teckenattribut (färg och understrykning) vars egenskaper hämtas från vissa teckenformatmallar.  
Om du inte vill ha den automatiska URL-igenkänningen finns det flera möjligheter att ta bort den:  
Ångra URL-igenkänning  
Om du håller på att skriva och en text just har omvandlats automatiskt till en hyperlänk kan du ångra den här formateringen genom att trycka på tangentkombinationen Kommando Ctrl +Z.  
Om du först senare märker att texten har omvandlats markerar du hyperlänken och väljer Format - Standard.  
Stänga av URL-igenkänning  
Ladda ett dokument av den typen som du vill ändra URL-igenkänningen för.  
Om du vill ändra URL-igenkänningen för textdokument öppnar du ett textdokument.  
Välj Verktyg - AutoKorrigering. (I %PRODUCTNAME Writer heter kommandot Verktyg - AutoKorrigering / AutoFormat.)  
I dialogrutan AutoKorrigering klickar du på fliken Alternativ.  
Om du avmarkerar Känn igen URL ersätts ord inte längre automatiskt med hyperlänkar.  
I %PRODUCTNAME Writer finns det två kryssrutor framför Känn igen URL: rutan i den första kolumnen gäller för senare redigering och rutan i den andra kolumnen gäller för AutoKorrigering under textinmatningen.  
Visa, dölja och förankra fönster  
Du kan dölja fönster som Gallery, Navigator och Stylist tillfälligt, i stället för att ständigt flytta eller öppna och stänga dem.  
Du kan välja om fönstren skall täcka det aktuella dokumentet eller om de delar utrymmet på bildskärmen med det aktuella dokumentet.  
Förankra fönster och göra dem till fria fönster  
Det finns två möjligheter:  
Håll ner Ctrl-tangenten och dra fönstret i titellisten till kanten.  
Håll ner Ctrl-tangenten och dubbelklicka på ett fritt område i fönstret eller på ett ställe i det gråa området i fönstret där ingen ikon finns.  
Men den här metoden kan du också göra ett förankrat fönster till ett fritt fönster igen.  
Visa och dölja förankrade fönster  
I kanten av ett förankrat fönster hittar du en kommandoknapp med en pin.  
Den används för att växla mellan "svävande" och "fixera ".  
Med den här kommandoknappen kan du välja om det förankrade fönstret visas tillsammans med det aktuella dokumentet eller om fönstret tillfälligt täcker dokumentet.  
Om du inte använder kommandoknappen med pilen för att visa fönstret utan bara klickar på den synliga kanten av det förankrade fönstret visas det inte permanent utan bara tillfälligt.  
Om du flyttar muspekaren en bit bort från ett fönster som visas tillfälligt, döljs det.  
AutoHide-funktionen arbetar oberoende av om du visar fönstret svävande eller fixerat.  
Om det är i fokus, när du alltså har klickat där, måste du klicka en gång utanför fönstret för att det skall döljas igen.  
Om fönstret inte är i fokus döljs det automatiskt.  
Beskrivningen i det här avsnittet gäller också för andra fönster som t.ex. Navigator, Stylist, Gallery eller förhandsvisningsfönstret i %PRODUCTNAME Impress.  
Om de här fönstren är förankrade och du sedan har visat dem genom att klicka på fönsterkanten för att använda AutoHide-funktionen, klickar du bara i det aktuella dokumentet och fönstret döljs.  
AutoHide-funktionen gäller alltid för alla fyra fönsterkanter för alla fönster som är förankrade i den här kanten.  
Definiera bakgrundsfärg eller bakgrundsgrafik  
Du kan definiera en bakgrundsfärg för olika objekt.  
Med en del objekt kan man t.o.m. ha ett grafikobjekt som bakgrund.  
Ge texttecken en bakgrund  
Markera tecknen.  
Välj Format - Tecken.  
Klicka på fliken Bakgrund och välj bakgrundsfärg.  
Ge stycke en bakgrund  
Placera markören i stycket eller markera flera stycken.  
Välj Format - Stycke.  
Klicka på fliken Bakgrund och välj en bakgrundsfärg eller ett bakgrundsgrafikobjekt.  
Förse texttabell helt eller delvis med bakgrund  
Placera markören i tabellen i ditt textdokument.  
Välj Format - Tabell.  
Klicka på fliken Bakgrund och välj en bakgrundsfärg eller ett bakgrundsgrafikobjekt.  
I ett fält väljer du om färgen eller grafikobjektet ska gälla för den aktuella cellen, den aktuella raden eller hela tabellen.  
Om du markerar flera celler eller rader innan du öppnar dialogrutan gäller ändringen för markeringen.  
Förse %PRODUCTNAME Calc-tabell med bakgrund  
Markera cellerna.  
Välj Format - Cell (eller Formatera celler på snabbmenyn).  
Klicka på fliken Bakgrund och välj en bakgrundsfärg.  
Grafik i bakgrunden till celler  
Välj Infoga - Grafik - Från fil.  
Välj ett grafikobjekt och klicka på Öppna.  
Grafikobjektet infogas i den aktuella cellen.  
Du kan flytta och skala grafikobjektet som du vill.  
På snabbmenyn hittar du kommandot Placering - I bakgrunden som du använder om du vill placera grafikobjektet i bakgrunden.  
Använd sedan Navigator Navigator om du vill markera grafikobjektet.  
Grafik i bakgrunden på utskrivna sidor (vattenmärke)  
Välj Format - Sida.  
Klicka på fliken Bakgrund och välj en bakgrundsfärg eller ett bakgrundsgrafikobjekt.  
Den här bakgrunden visas bara på utskrift bakom de celler som inte annars är formaterade.  
Ge presentationssidor en bakgrund  
Se.  
Fliken Bakgrund  
Definiera inramning  
Du kan definiera inramningar av sidor, tabeller och andra objekt på två ställen:  
Meny Format - (Objektnamn) - Inramning  
Utrullningslist Inramning på objektlisten när objektet är markerat (gäller inte för alla objekt).  
Meny Format, använd fliken Inramning  
Använd utrullningslisten Inramning  
Anta att du vill använda följande tabellinramning i ett dokument:  
1.  
Ställ markören på det ställe i dokumentet där tabellen ska infogas.  
2.  
Öppna dialogrutan Infoga tabell med menykommandot Infoga - Tabell och infoga en tabell med önskad storlek, t.ex. 3 kolumner och 5 rader.  
3.  
Markera hela tabellen, tryck på tangentkombinationen Ctrl+A två gånger, och klicka på ikonen Inramning.  
På utrullningslisten klickar du på ikonen som finns uppe till vänster och som symboliserar "Ingen inramning".  
4.  
Markera nu hela den första raden med musen och öppna dialogrutan Tabellformat med snabbmenykommandot Tabell.  
5.  
Klicka på fliken Inramning.  
6.  
Välj linjetjocklek i fältet Linje, t.ex. 2,50 pt.  
7.  
Klicka en gång på området mellan de båda undre vinklarna (se illustration) i det stora fältet Linjeplacering och sedan på OK.  
8.  
Markera nu kolumnen i mitten av tabellen och öppna dialogrutan Tabellformat igen via snabbmenykommandot Tabell.  
9.  
Klicka på områdena som representerar den högra och vänstra linjen under Linjeplacering, se illustration.  
10.  
Definiera linjetjockleken i fältet Linje och klicka på OK.  
11.  
Markera den understa raden i tabellen och öppna dialogrutan Tabellformat igen via snabbmenykommandot Tabell.  
12.  
Välj linjetjocklek i fältet Linje, hittills 2,50 pt, och klicka sedan på områdena som representerar den övre och undre linjen under Linjeplacering.  
13.  
Klicka sedan på OK så är tabellen färdig.  
Fliken Inramning  
Ändra rubrik på ett dokument  
På titellisten visar %PRODUCTNAME bl.a. rubriken på det aktuella dokumentet.  
Om du skapar och sparar ett nytt dokument är rubriken identisk med filnamnet.  
Så här ändrar du rubriken på det aktuella dokumentet  
Välj Arkiv - Egenskaper.  
Dialogrutan Egenskaper för öppnas.  
Klicka på fliken Beskrivning.  
Mata in rubriken i textfältet Rubrik och klicka på OK.  
Egenskaper för  
Redigera diagramaxel  
Anta att du har infogat ett diagram i t.ex. ett %PRODUCTNAME Calc-dokument och vill ändra skalan för den lodräta Y-axeln.  
Dubbelklicka på diagrammet.  
Diagrammet får gråa kanter och menylisten visar nu kommandon för redigering av objekt i diagrammet.  
Välj Format - Axel - Y-axel om du vill redigera Y-axeln eller dubbelklicka på Y-axeln.  
Dialogrutan Y-axel öppnas.  
Klicka t.ex. på fliken Skalning om du vill ändra axelns skala.  
Klicka på OK.  
I ditt dokument klickar du utanför diagrammet för att lämna redigeringsläget för diagrammet.  
Format - Objektegenskaper  
Förse diagramstaplar med textur  
Tilldela en stapeltyp en bitmap (i stället för t.ex. en opak färg):  
Växla till redigeringsläget genom att dubbelklicka på diagrammet.  
Dubbelklicka på motsvarande stapel (alla staplar med den här färgen är nu markerade).  
Välj Objektegenskaper på snabbmenyn, sedan fliken Yta.  
Klicka på Bitmap.  
I listrutan kan du nu välja ut en bitmap som textur för den här stapeln.  
Genom att klicka på OK övertar du inställningen.  
AutoPilot Diagram  
Infoga diagram  
1.  
Öppna ett tabelldokument och skriv lite data med rad - och kolumnrubriker i en tabell.  
2.  
Markera uppgifterna tillsammans med överskrifterna.  
3.  
Klicka på ikonen Infoga diagram på utrullningslisten Infoga objekt på verktygslisten.  
Markören blir till ett hårkors med en diagramsymbol.  
4.  
I tabelldokumentet ritar du upp en rektangel som anger platsen och storleken för diagrammet.  
Båda går att ändra i efterhand.  
När du släpper musknappen öppnas en dialogruta där du kan göra fler inmatningar eller klicka på kommandoknappen Färdigställ för att skapa diagrammet med standardinställningarna.  
Vi visar här ett exempel (dokument Bio1.sxc i exempelmappen) där du kan se antalet biobesökare i olika åldersgrupper för olika städer.  
Om du hellre vill ha städerna på den horisontella axeln i stället för åldersgrupperna, kan du "tippa" diagrammet i efterhand.  
Så länge diagrammet är markerat hittar du ikonen Data i kolumner på verktygslisten.  
Klicka på den!  
Det är möjligt att göra fler ändringar av de enskilda elementen i diagrammet.  
Du kan antingen dubbelklicka på de enskilda delarna i diagrammet eller välja de enskilda alternativen på menyn Format vid aktiverat diagram.  
Om du till exempel dubbelklickar på färgförhandsvisningen i förklaringen så kan du automatiskt formatera alla tillhörande datapunkter på nytt.  
Om du däremot klickar på bakgrunden i rutan med förklaringen så formaterar du bakgrunden till förklaringen.  
Om du har skapat diagrammet med data från en %PRODUCTNAME Calc-tabell markeras dataserierna i tabellen när du klickar på dem i diagrammet.  
Du kanske har ställt diagrammet i din %PRODUCTNAME Calc-tabell i bakgrunden och undrar nu hur du kan markera det för vidare redigering?  
Öppna utrullningslisten Visa ritfunktioner och välj det första verktyget, Urval spilen.  
Med den kan du klicka på diagrammet.  
Det är möjligt att flytta en dataserie framåt eller bakåt i ett diagram i %PRODUCTNAME Calc.  
Du kan placera serierna på ett sådant sätt så att de lägsta 3D-visningarna står längst fram och de högre längre bak.  
För att ändra placeringen i diagrammet använder du ett kommando på snabbmenyn till en dataserie resp. under Format - Placering.  
Utgångsdata i %PRODUCTNAME Calc-tabellen placeras inte om.  
Om du infogar ett diagram via utrullningslisten Infoga - Infoga diagram i ett presentations - eller teckningsdokument visas det med en uppsättning av exempeldata.  
Om du vill infoga ett diagram i ett tabelldokument måste du markera cellerna i tabellen vars värden skall visas i diagrammet.  
Även i ett %PRODUCTNAME Writer-dokument kan du infoga ett diagram som bygger på data från en %PRODUCTNAME Writer-tabell.  
Om du inte har markerat några data i en %PRODUCTNAME Writer-tabell infogar menykommandot Infoga - Objekt - Diagram ett diagram med exempeldata även i %PRODUCTNAME Writer.  
Du kan ändra värdena i ett diagram med exempeldata genom att dubbelklicka på diagrammet och sedan välja Redigera - Diagramdata.  
Om du vill ändra värdena i ett diagram som bygger på markerade data, måste du ändra värdena i tabellens celler.  
Om det rör sig om ett diagram i ett textdokument, trycker du på F9 för att uppdatera diagrammet.  
Du har också möjlighet att ändra diagramdata om du har kopierat ett diagram från t.ex. ett %PRODUCTNAME Calc-dokument till ett %PRODUCTNAME Writer-dokument och sedan dubbelklickar på det i %PRODUCTNAME Writer-dokumentet.  
Men då redigerar du bara en kopia som inte har någon förbindelse till de ursprungliga värdena i tabellen.  
Du kan ändra diagramtypen i efterhand.  
I dialogrutan som öppnas när du har dubbelklickat på diagrammet och valt Format - Diagramtyp kan du välja bland de olika typerna.  
Växla också mellan 2D - och 3D-visningarna.  
Vid typen Staplar kan du välja Kombinationsdiagram av staplar och linjer.  
De tredimensionella visningarna gör att det är möjligt att använda särskilda effekter.  
För 3D-diagram kan du till och med ställa in belysning, omgivningsljus och färgfilter.  
3D-diagram kan du rotera och tippa interaktivt med musen för att justera dem optimalt.  
XY-diagram kan du förse med statistiska värden via kommandot Infoga - Statistik, t.ex. felindikatorer för varians, med regressionskurvor och mycket annat.  
Även en enkel eller dubbel logaritmisk visning av axlarna går att ställa in här.  
I linjediagram kan du arbeta med olika symboler som du antingen kan låta %PRODUCTNAME sätta in automatiskt eller välja ut från grafikfiler eller Gallery.  
AutoPilot Diagram  
Redigera diagramförklaring  
Anta att du har infogat ett diagram i t.ex. ett %PRODUCTNAME Calc-dokument och vill ge förklaringen en färggradient.  
Dubbelklicka på diagrammet.  
Diagrammet får gråa kanter och menylisten visar nu kommandon för redigering av objekt i diagrammet.  
Välj Format - Förklaring eller dubbelklicka på förklaringen.  
Dialogrutan Förklaring öppnas.  
Klicka t.ex. på fliken Yta om du vill ändra förklaringens bakgrund.  
Välj Färggradient i kombinationsfältet och välj en färggradient på listan.  
Klicka på OK.  
I ditt dokument klickar du utanför diagrammet för att lämna redigeringsläget för diagrammet.  
I %PRODUCTNAME Draw definierar du egna färggradienter, skrafferingar, bitmaps och färger.  
Om du vill markera förklaringen dubbelklickar du först på diagrammet (se steg 1) och klickar sedan på förklaringen.  
Du kan nu flytta förklaringen inuti diagrammet med musen.  
Om du har flyttat förklaringen över ett annat objekt i diagrammet kan du inte längre öppna förklaringens egenskapsdialog genom att dubbelklicka.  
När du vill öppna egenskapsdialogen använder du antingen menyn Format eller klickar en gång på förklaringen och sedan öppnar du snabbmenyn och väljer Objektegenskaper.  
Motsvarande gäller för alla andra objekt i diagrammet.  
Format - Objektegenskaper  
Redigera diagramrubrik  
Anta att du har infogat ett diagram i t.ex. ett %PRODUCTNAME Calc-dokument och vill ändra rubriken.  
Dubbelklicka på diagrammet.  
Diagrammet får gråa kanter och menylisten visar nu kommandon för redigering av objekt i diagram.  
Dubbelklicka på standardrubriktexten.  
Texten får en grå kant och du kan ändra den.  
Med returtangenten skapar du en ny rad.  
Om du klickar enkelt på rubriken i stället för att dubbelklicka kan du flytta den med musen.  
Välj Format - Rubrik - Huvudrubrik om du vill redigera formateringen av huvudrubriken.  
Dialogrutan Rubrik öppnas.  
Klicka t.ex. på fliken Tecken om du vill ändra teckensnittet.  
Klicka på OK.  
I ditt dokument klickar du utanför diagrammet för att lämna redigeringsläget för diagrammet.  
Format - Objektegenskaper  
Anpassa tangentbord  
Du kan lägga till alla okända ord som finns i ett textdokument i den aktiverade användarordlistan med ett enda kommando.  
Men du måste själv lägga kommandot på en tangentkombination eller en ikon först.  
Öppna ett valfritt textdokument.  
Välj Verktyg - Anpassa...  
Dialogrutan Anpassa visas.  
Om du vill tilldela en tangentkombination klickar du på fliken Tangentbord.  
Om du vill lägga till en egen ikon för den här funktionen på en symbollist klickar du på fliken Symbollister.  
Här beskriver vi hur du anpassar tangentkombinationer.  
Hur du placerar en ny ikon på en symbollist beskrivs under Skapa en faxikon.  
Markera sedan Lägg till okända ord i listrutan Funktion.  
Sök nu i den stora listrutan Tangentkombinationer efter en ledig tangentkombination för det här kommandot (t.ex. F10).  
Klicka på Ändra och stäng dialogrutan med OK.  
Genom att trycka på den tangent eller tangentkombination som du har valt kan du nu göra så att en rättstavningskontroll genomförs i det aktuella textdokumentet och att alla okända ord automatiskt läggs till i en aktiverad användarordlista.  
Följande villkor måste uppfyllas för att de okända orden ska kunna läggas till:  
Användarordlistan ska vara aktiverad.  
Användarordlistan får inte vara någon negativ-ordlista.  
Språket i användarordlistan måste vara inställd på "alla".  
Användarordlistans fil får inte vara skrivskyddad.  
Verktyg - Anpassa  
Anpassa meny  
För att du ska kunna integrera en skanner krävs en lämplig skannerdrivrutin som passar ditt operativsystem.  
För tillfället kan TWAIN-drivrutiner i Windows och SANE-drivrutiner i Unix integreras i %PRODUCTNAME.  
Det exempel som visas här för att integrera kommandon på en %PRODUCTNAME -meny kan också användas för andra funktioner, oberoende av om det rör sig om en skanner eller inte.  
I modulerna för redigering av grafik har %PRODUCTNAME även menykommandon för skanning.  
Dessa fungerar om du har integrerat en TWAIN-kompatibel drivrutin för din skanner eller din digitala kamera i systemet.  
Här beskrivs hur du integrerar skanningskommandon på Arkivmenyn i ett textdokument.  
En TWAIN-drivrutin infogas för det mesta på arkivmenyn.  
Där ska vi lägga in posten "Skanna", som i sin tur ska ha de två underordnade posterna "Välj källa" och "Skanna in ".  
De respektive dialogrutorna och funktionerna som aktiveras och utförs när dessa poster har valts kommer från TWAIN-drivrutinen. %PRODUCTNAME anropar dem bara.  
Öppna ett textdokument som aktivt dokument.  
Välj Verktyg - Anpassa....  
Dialogrutan Anpassa visas.  
Klicka på fliken Meny.  
I den stora listrutan klickar du på det kommando under vilket du vill placera skanningskommandot, t.ex. på "Versioner".  
Klicka på kommandoknappen Ny meny.  
Under den senast markerade posten ser du en ny post med namnet "Meny".  
Den har redan en underordnad post som är en skiljelinje.  
Klicka två gånger efter varandra med höger musknapp på den nya posten "Meny" och mata in det nya namnet "Skanna ".  
Klicka på den underordnade posten, d.v.s. linjen.  
Om du nu definierar nya menyposter förs dessa in som undermenyer till "Skanna".  
I den vänstra listrutan väljer du funktionskategorin "Infoga" och sedan i höger listruta funktionen "Skanningskälla ".  
Det nya menykommandot infogas i den stora listrutan.  
Välj funktionen "Beställ en skanning" i den högra listrutan och klicka återigen på Nytt.  
Även den här posten fogas in.  
Klicka på skiljelinjen och sedan på Radera.  
Strecket tas bort.  
Om du vill kan du också döpa om de båda undermenyposterna (klicka på dem med höger musknapp).  
Genom att dra och släppa flyttar du om namnen i den stora listrutan.  
Ändringarna sparas automatiskt.  
Från och med nu har du alltid tillgång till de nya menyposterna.  
Verktyg - Anpassa  
Anpassa %PRODUCTNAME  
Du kan skräddarsy %PRODUCTNAME.  
Posterna på menylisten kan du redigera hur du vill: du kan radera poster, lägga till nya, kopiera eller flytta poster från en meny till en annan, byta namn på dem och så vidare.  
Du kan konfigurera symbollisterna som du vill.  
Ikoner kan du flytta genom att hålla ner Alt-tangenten och använda dra-och-släpp (i Windows).  
Du kan ändra tangentkombinationer efter dina önskemål.  
Du gör sådana ändringar i dialogrutan som öppnas via Verktyg - Anpassa.  
Verktyg - Anpassa  
Spara konfiguration med ett dokument  
Du kan om du vill definiera en konfiguration globalt (då gäller den alltid när du senare aktiverar ett dokument av samma typ som när du definierade konfigurationen), eller också kan du koppla en konfiguration till ett visst dokument, som i så fall måste finnas som fil när du gör det.  
Ladda det dokument som du vill koppla konfigurationen till, eller aktivera ett valfritt dokument av samma typ.  
Ställ in konfigurationen.  
Välj t.ex. vilka symbollister som ska vara synliga, eller definiera innehållet på symbollisterna, posterna på menyerna eller på statuslisten och så vidare.  
Alla inställningsmöjligheter finns sammanfattade i dialogrutan Verktyg - Anpassa...  
Klicka på kommandoknappen Spara... i dialogrutan Verktyg - Anpassa...  
Dialogrutan för att spara konfigurationen visas.  
I listrutan Filtyp väljer du <Alla>.  
I den stora listrutan i dialogrutan Spara väljer du sedan den fil som du vill koppla konfigurationen till.  
Klicka på Spara...  
Du får nu en fråga om du vill ersätta den aktuella filen.  
Den frågan gäller i det här fallet bara den konfiguration som eventuellt redan är kopplad till dokumentet och inte dokumentets "egentliga" innehåll.  
Bekräfta därför överskrivningen.  
Nu är den aktuella konfigurationen kopplad till det valda dokumentet.  
Du kan kontrollera detta genom att ladda dokumentet, öppna dialogrutan Arkiv - Dokumentmall - Administrera och där dubbelklicka på dokumentet.  
Varje gång som du laddar eller aktiverar dokumentet, aktiveras också den konfiguration som har sparats tillsammans med det.  
Om du aktiverar eller laddar ett annat dokument, som inte innehåller någon konfigurationsinformation, används återigen den globala standardkonfigurationen.  
Denna kan du alltid ställa in för hand genom att öppna dialogrutan Verktyg - Anpassa... och klicka på kommandoknappen Återställ.  
Verktyg - Anpassa  
Kopiera ritobjekt till ett annat dokument  
I %PRODUCTNAME går det att kopiera ritobjekt direkt mellan text - tabell - och presentationsdokument.  
Markera ett eller flera ritobjekt.  
Kopiera ritobjektet till urklippet genom att t.ex. trycka på Kommando Ctrl +C.  
Växla till det andra dokumentet och placera markören där ritobjektet ska klistras in.  
Klistra in ritobjektet, t.ex. genom att trycka på Kommando Ctrl +V.  
Klistra in i ett textdokument  
Ett inklistrat ritobjekt är förankrat i det aktuella stycket i ett textdokument.  
Du kan byta förankring genom att markera objektet och klicka på ikonen Byt förankring på objektlisten.  
En popupmeny öppnas där du kan välja mellan olika typer av förankring.  
Klistra in i ett tabelldokument  
Ett inklistrat ritobjekt är förankrat i den aktuella cellen i ett tabelldokument.  
Du kan byta förankring mellan cell och sida och tillbaka genom att markera objektet och klicka på ikonen Byt förankring.  
Klistra in data från tabelldokument  
Om du bara vill kopiera innehållet (text eller siffror) i en cell gör du detta via urklippet.  
Även formlerna som står i cellerna kan kopieras från formellistens inmatningsrad till urklippet och sedan klistras in i en text.  
Använd sedan urklippet eller dra-och-släpp och klistra in cellerna i textdokumentet.  
I textdokumentet hittar du sedan ett OLE-objekt som du kan fortsätta att redigera som du vill.  
Om du drar tabellcellerna till teckningsvyn i ett presentationsdokument placeras de som OLE-objekt även där.  
Varje tabellcell utgör en rad i dispositionsvyn.  
Cellerna flyttas när du använder dra-och-släpp.  
Det är bara om du håller ner skifttangenten när du drar som de kopieras.  
Klistra in data från textdokument  
Du kan överföra texter till andra dokumenttyper som tabelldokument och presentationer.  
Du måste välja om texten ska sättas i en egen textram eller placeras i en tabellcell eller i dispositionen till en presentation.  
Om du överför texten via urklippet kan du klistra in den igen med eller utan textattribut på önskat ställe.  
Använd tangentkombinationerna för Kopiera Kommando Ctrl +C och Klistra in Kommando Ctrl +V.  
För att välja formatet med vilket urklippets innehåll ska klistras in, klickar du lite längre på ikonen Klistra in på funktionslisten.  
På undermenyn väljer du ut ett format.  
Ett motsvarande urval av format finns under Redigera - Klistra in innehåll.  
Om du utgår från ett textdokument finns kommandot Skicka - Disposition till presentation på Arkiv -menyn.  
Ett nytt presentationsdokument skapas där överskrifterna från textdokumentet utgör dispositionen.  
Det här kommandot visas bara om överskrifterna är formaterade med en motsvarande styckeformatmall.  
Om du även vill använda det första underordnade stycket (eller flera stycken) från texten väljer du AutoUtdrag till presentation.  
Det här kommandot visas bara om överskrifterna är formaterade med en motsvarande styckeformatmall.  
Kopiera text med dra-och-släpp  
Om du markerar ett textavsnitt och sedan drar det till ett tabelldokument infogas det som text i den cell där du släpper musknappen.  
Om du drar ett textavsnitt till teckningsvyn i ett presentationsdokument infogas ett OLE-objekt som %PRODUCTNAME -plug-in.  
Om du drar texten till dispositionsvyn i en presentation infogas den vid markören.  
Registrera adressbok  
I %PRODUCTNAME kan du registrera olika datakällor.  
Innehållet i datafälten är då tillgängliga i t.ex. fältkommandon och kontrollfält.  
Adressboken, som du kanske redan använder i ditt system, är en sådan datakälla, t.ex. en LDAP-server eller en Netscape-adressbok.  
I mallarna och AutoPiloterna i %PRODUCTNAME används fältkommandon för innehållet i adressboken.  
Eftersom det är omöjligt att veta vilken adressbok du använder i ditt system används först allmänna fältkommandon i mallarna.  
De allmänna fältkommandona fylls automatiskt med konkreta fältkommandon som är relevanta för ditt system första gången mallarna öppnas.  
För att den här ersättningen ska fungera måste du meddela %PRODUCTNAME vilken adressbok du använder.  
Dialogrutan där du gör det startar automatiskt när du t.ex. öppnar en mall till ett affärsbrev första gången.  
Du kan också öppna dialogrutan så här:  
AutoPilot för adressdatakällor  
Den här AutoPiloten öppnar du genom att välja Arkiv - AutoPilot - Adressdatakälla.  
Den beskrivs i %PRODUCTNAME -hjälpen.  
Registrera en adressbok manuellt  
1.  
Välj Arkiv - Dokumentmall - Adressbokskälla.  
Dialogrutan Mallar: adressbokstilldelning öppnas.  
2.  
Välj systemadressboken i fältet Datakälla eller datakällan som du vill använda som adressbok.  
Om du inte har registrerat systemadressboken som datakälla i %PRODUCTNAME än, klickar du på Administrera.  
Du kommer då till dialogrutan Administrera datakällor där du registrerar din systemadressbok som en ny datakälla i %PRODUCTNAME.  
Under Systemadressbok som datakälla nedan kan du läsa om hur du gör.  
3.  
I fältet Tabell väljer du databastabellen som du vill använda som adressbok.  
4.  
I området Fälttilldelning kan du nu definiera hur de fördefinierade fältnamnen för företag, avdelning, förnamn, efternamn och så vidare ska användas på de konkreta namnen i din adressbok.  
För en datakälla på engelska skulle du t.ex. öppna fältet bredvid posten Företag och där t.ex. välja ut Company.  
I fältet bredvid Avdelning väljer du Department och så vidare.  
Stäng dialogrutan med OK.  
5.  
Från och med nu är din datakälla känd som adressbok i %PRODUCTNAME.  
Om du öppnar en mall från kategorin Affärskorrespondens kan %PRODUCTNAME automatiskt använda fältkommandona för ett standardbrev (kopplad utskrift) på rätt sätt.  
Systemadressbok som datakälla  
1.  
Dialogrutan Administrera datakällor öppnas om du väljer Arkiv - Dokumentmall - Adressbokskälla och klickar på Administrera (se anvisningar ovan) eller om du väljer Verktyg - Datakällor.  
2.  
Klicka på kommandoknappen Ny datakälla.  
3.  
Välj Adressbok under Databastyp.  
4.  
Klicka på... för att öppna dialogrutan Datakälla.  
5.  
Välj datakälla och klicka på OK.  
Om du har valt LDAP adressbok har nu dialogrutan Administrera datakällor en ny flik som heter LDAP där du kan ange LDAP-servern och dess parametrar.  
6.  
Klicka på fliken Tabeller.  
Markera tabellerna som ska visas i %PRODUCTNAME.  
7.  
Under fliken Allmänt kan du ange ett namn för den här datakällan i fältet Namn.  
Stäng dialogrutan med OK.  
Administrera datakällor  
Datakällöversikt  
Datakällvy  
Du öppnar datakällvyn med Visa - Datakällor (F4) från ett text - eller tabelldokument.  
Till vänster ser du Explorer för datakällor.  
Om du markerar en tabell eller sökning där visas innehållet i tabellen eller sökningen till höger.  
I övre kanten finns Databaslisten.  
Datakällor  
Registrera ny datakälla, Adressbok som datakälla  
Redigera datakällnamn eller typ  
Titta på innehåll i datakällor  
Tabeller  
Skapa nu tabell, redigera struktur, Index, Relationer  
Mata in, redigera och kopiera dataposter  
Sökningar  
Skapa ny sökning, redigera struktur  
Mata in, redigera och kopiera dataposter  
Formulär  
Skapa nya formulädokument, Redigera formulärfunktioner  
Titta på formulärdokument, Mata in resp. redigera formulär  
Övrigt  
Snabbmenyer i Explorer för datakällor (till vänster)  
Snabbmenyer i datakällvyn (till höger  
Import och export av data i textformat  
Om du vill utbyta data med en databas, som inte har en ODBC-koppling och inte tillåter någon dBase-import och -export, så kan du oftast utbyta data genom att använda ett gemensamt textformat.  
Import av data till %PRODUCTNAME  
För utbyte av data i textformat använder du import - och exportfiltren från %PRODUCTNAME Calc:  
Exportera önskade data från källdatabasen i ett textformat.  
Det är bäst att välja CSV-textformat, där datafälten t.ex. är avskilda med komman och dataposterna med radbrytningar.  
Öppna dessa data med hjälp av filfiltret "Text CSV".  
Du väljer det här filfiltret i dialogrutan Öppna i listrutan Filtyp.  
Välj filen och bekräfta med Öppna.  
Du ser dialogrutan Textimport.  
Här kan du i stor utsträckning ställa in vilka data du vill använda från textdokumentet.  
Så snart du har tillgång till dessa data i en %PRODUCTNAME Calc-tabell, kan du redigera dem.  
Det finns två sätt att spara data i en %PRODUCTNAME -datakälla.  
Spara den aktuella %PRODUCTNAME Calc-tabellen i dBase-format i mappen till en dBase-databas.  
För att göra detta väljer du Arkiv - Spara som, sedan väljer du Filtyp "dBase" och mappen för dBase-databasen.  
Markera dataområdet i %PRODUCTNAME Calc-tabellen och dra området till en tabellcontainer i datakällvyn.  
Tabellcontainern är området med beteckningen "Tabeller" till vänster i databas-Explorer (se bild).  
En AutoPilot startas automatiskt.  
Export till csv-textformat  
Den aktuella %PRODUCTNAME -tabellen kan du exportera i ett textformat som kan läsas av många andra program.  
Välj Arkiv - Spara som.  
I fältet Filtyp väljer du filtret "Text CSV".  
Mata in ett filnamn och klicka på Spara.  
Dialogrutan Textexport öppnas där du kan välja teckenuppsättning, fältavgränsare och textavgränsare.  
Klicka på OK.  
Du får information om att bara den aktuella tabellen har sparats.  
Utföra SQL-kommando direkt  
Det går även att styra en databas direkt med hjälp av SQL-kommandon, skapa, redigera tabeller, skapa sökningar och så vidare.  
Det går inte att använda alla SQL-anvisningar i alla databastyper.  
Ta reda på vilka SQL-kommandon som understöds av ditt databassystem.  
1.  
Öppna dialogrutan Administrera datakällor via Verktyg - Datakällor.  
2.  
I listan markerar du datakällan som du vill anropa direkt via SQL och välj sidan Sökningar.  
3.  
Klicka på ikonen Mata in nytt SQL-kommando eller  
välj en befintlig sökning från listan och klicka på ikonen Mata in SQL-kommando.  
4.  
I dialogrutan Sökning matar du in SQL-kommandot som du vill utföra eller ändrar ett befintligt kommando enligt dina krav.  
5.  
Klicka på ikonen Utför.  
Resultatet av sökningen visas i det övre fönstret.  
6.  
Klicka på ikonen Spara eller Spara som för att spara den skapade eller ändrade sökningen.  
Ladda data från datakällor i %PRODUCTNAME Calc  
Om du bara vill exportera några dataposter från en datakälltabell markerar du dataposterna genom att klicka på radhuvudena.  
Använd skifttangenten och / eller Kommando Ctrl -tangenten för att göra en multimarkering.  
Släpp inte musknappen när du har markerat den sista dataposten utan dra de markerade dataposterna med nedtryckt musknapp till en öppen %PRODUCTNAME Calc-tabell.  
Nu kan du spara %PRODUCTNAME Calc-tabellen i ett valfritt format.  
Söka med ett formulärfilter  
1.  
Öppna ett formulär.  
Stäng av utkastläget.  
För att snabbt prova funktionen:  
Öppna ett tomt textdokument, tryck på F4, öppna litteraturdatabastabellen biblio i datakällvyn.  
Håll ner Skift+Ctrl-tangenterna och dra några kolumnhuvuden till dokumentet så att formulärfält skapas där.  
2.  
Stäng av utkastläget.  
För att göra det öppnar du utrullningslisten Formulärfunktioner och klickar på ikonen Utkastläge på / av så att den inte är intryckt.  
3.  
På formulärlisten klickar du på ikonen Formulärbaserat filter.  
Det aktuella formuläret visas med sina infogade formulärfunktioner som tom inmatningsmask.  
Vid den undre kanten visas Filterlisten.  
4.  
Du anger filtervillkoren i ett eller flera fält.  
Information om platshållare och operatorer som du kan använda finns i hjälpen för sökningsutkast.  
Om du anger filtervillkor i flera fält, kopplas de ihop med den logiska operatorn OCH.  
Om du klickar på ikonen Använd filter på filterlisten, utförs filtreringen i databasen.  
Formulärlisten visas igen och du kan navigera mellan träffarna.  
Om du klickar på kommandoknappen Stäng på filterlisten, visas formuläret utan filter.  
I formulärvyn kan du växla till filtrerad vy med ikonen Använd filter.  
Du kan ta bort det satta filtret med ikonen Ta bort filter / sortering.  
Om du vill koppla ihop flera filtervillkor med ELLER, klickar du på ikonen Filternavigation på filterlisten.  
Då öppnas det förankringsbara fönstret Filternavigator.  
När du sätter ett filter visas en tom filternivå längst ner i Filternavigator.  
Så snart du har markerat den kan du mata in fler filtervillkor i formuläret.  
Villkoren kopplas ihop med de redan inmatade med ett logiskt ELLER.  
För varje post i Filternavigator kan du öppna en snabbmeny.  
Här kan du direkt redigera filtervillkoren som text.  
Dessutom kan du välja filtervillkoren "Är tom" (SQL:  
Is Null) eller "Är inte tom "(SQL:  
Is not Null) om du vill undersöka om ett fält har något innehåll eller ej.  
Via snabbmenyn kan du också radera en post.  
Om du samtidigt håller ned Kommando Ctrl -tangenten kopieras de.  
Söka i tabeller och formulärdokument  
I tabeller och dokument där formulärfunktioner används, kan du öppna en dialogruta genom att klicka på ikonen Sök datapost med vars hjälp du kan hitta valfria texter och värden.  
Använd ikonen nere på formulärlisten, inte ikonen med liknande utseende på den vänstra verktygslisten.  
Du kan söka i ett bestämt datafält i alla dataposter eller i alla datafält.  
Du kan välja om texten ska stå i början av ett datafält, i slutet eller var som helst i fältet.  
Dessutom kan du arbeta med jokertecknen? och * eller med reguljära uttryck som i dialogrutan Sök och ersätt.  
I %PRODUCTNAME -hjälpen finns det mer information om sökfunktionen för databaser.  
Tabellutkast  
Här ser du hur du skapar en ny databastabell i utkastvyn.  
Öppna datakällvyn (F4).  
Där öppnar du en datakälla genom att klicka på plustecknet framför namnet.  
Tabellcontainern som kallas "Tabeller" visas.  
Nu öppnar du snabbmenyn genom att högerklicka på tabellnamnet.  
Skapa en ny tabell genom att välja Nytt tabellutkast.  
Du kan nu definiera datafälten i utkastvyn.  
Nya datafält matar du in rad för rad uppifrån och ned.  
För varje nytt datafält klickar du i cellen längst till vänster och anger ett fältnamn.  
I nästa cell till höger bestämmer du fälttyp.  
När du klickar i cellen visas en listruta där du kan välja mellan olika fälttyper.  
Varje enskilt datafält kan bara innehålla data som motsvarar den fälttyp som du har definierat.  
Du kan t.ex. inte mata in text i ett talfält.  
I dem kan du mata in upp till 64 kB text.  
Du kan även göra en beskrivning till varje datafält.  
Beskrivningens text visas i tipshjälpen för kolumnhuvudena i tabellvyn.  
Fältegenskaper  
Här matar du in egenskaper för varje markerat datafält.  
Vilka inmatningsmöjligheter som är tillgängliga beror på databastypen.  
Under Standardvärde ger du datafältet ett innehåll som ska finnas i alla nya dataposter, men som naturligtvis går att ändra.  
Under Inmatning krävs anger du om datafältet får vara tomt eller inte.  
Vilka urvalsmöjligheter som är tillgängliga i listrutan för Fältlängd beror på vald fälttyp.  
Det är bara utkastvyn som får vara öppen.  
Spara dokument automatiskt  
Spara en säkerhetskopia varje gång du sparar  
Öppna dialogrutan Verktyg - Alternativ - Ladda / spara - Allmänt.  
Markera rutan Skapa alltid säkerhetskopia.  
Om du sparar det aktuella dokumentet med Arkiv - Spara eller Ctrl+S och använder filnamnet och sökvägen som du har öppnat dokumentet ifrån, skrivs den gamla versionen över av den nya.  
Om rutan Skapa alltid säkerhetskopia är markerad kopieras den gamla versionen först till Backup-katalogen.  
Backup-katalogen heter {installpath} / user / backup {installpath }\user\backup.  
Du kan ändra den i dialogrutan Verktyg - Alternativ - %PRODUCTNAME - Sökvägar vid "Säkerhetskopior".  
Kopian har samma namn som dokumentet men filtillägget .BAK.  
Om det redan finns en fil med det namnet i Backup-katalogen, skrivs den över utan kontrollfråga!  
Spara automatiskt var n minut  
Öppna dialogrutan Verktyg - Alternativ - Ladda / spara - Allmänt.  
Markera rutan Spara automatiskt var och välj tidsintervall i rotationsfältet.  
I dialogrutan kan du bestämma om du vill spara eller inte.  
Det här kommandot sparar det aktuella dokumentet, som om du t.ex. hade tryckt på Ctrl+S.  
Om dokumentet redan har sparats innan skrivs den gamla versionen över av den aktuella!  
Om du har aktiverat både Skapa alltid säkerhetskopia och Spara automatiskt var, skrivs filen över var n minut och samtidigt ersätts säkerhetskopian med den senaste versionen.  
Spara som  
Verktyg - Alternativ - Ladda / spara - Allmänt  
Öppna dokument  
Öppna ett existerande dokument  
Tryck på tangentkombinationen Kommando Ctrl +O.  
Dialogrutan Öppna visas.  
Välj en fil och klicka på Öppna.  
När du ska byta enhet anger du bara enhetsbokstaven med efterföljande kolon i textfältet Filnamn, t.ex. "c:" och trycker på returtangenten.  
Sedan visas direkt innehållet på C: i urvalsfönstret.  
Även i textfältet Filnamn i dialogrutan Öppna kan du skriva in en URL, som dock i helt utskriven form måste börja med file: / / / eller ftp: / / eller http: / /.  
Begränsa visningen av namn i Öppna-dialogrutan  
Vill du bara välja en av teckningarna bland alla dokumenten i en katalog?  
Välj Filtyp i fältet med samma namn i dialogrutan Öppna.  
Filtyperna är indelade i grupper.  
Om du t.ex. väljer posten Teckningar visas bara teckningsdokumenten som %PRODUCTNAME kan öppna i dialogrutan. %PRODUCTNAME bedömer detta efter filnamnstilläggen.  
Öppna dokument med samma sidposition (t.ex. på sidan 30) som det stängdes med  
Markera rutan Redigeringsvy under Verktyg - Alternativ - %PRODUCTNAME - Vy.  
Öppna ett tomt dokument  
Det finns flera möjligheter att öppna ett tomt dokument.  
Detta är en av dem:  
Klicka kort på ikonen Nytt på funktionslisten.  
Då öppnas ett dokument av den dokumenttyp som visas på ikonen.  
Om du håller ner musknappen lite längre på ikonen Nytt öppnas en undermeny där du kan välja en annan dokumenttyp.  
Arkiv - Öppna  
Spara dokument  
Tryck på tangentkombinationen Kommando Ctrl +S.  
Dokumentet arkiveras med sin sökväg och sitt namn på det aktuella lokala datamediet, nätverksenheten eller på Internet och skriver över en eventuell gammal version som kan finnas där.  
När du sparar en fil för första gången, visas dialogrutan Spara som där kan ange namn, katalog och enhet resp. volym för filen.  
Du öppnar den här dialogrutan via menykommandot Arkiv - Spara som.  
Du kan göra inställningar som t.ex. spara automatiskt eller skapa säkerhetskopia automatiskt under Verktyg - Alternativ - Ladda / spara - Allmänt.  
Spara som  
Verktyg - Alternativ - Ladda / spara - Allmänt  
Dra-och-släpp med datakällvy  
Det enklaste och snabbaste sättet att överföra data från en datakälla till ett text - eller tabelldokument, eller skapa formulär baserade på en datakälla, är dra-och-släpp-metoden.  
Kopiera med dra-och-släpp  
Om du har gjort fel vid dra-och-släpp och vill återställa funktionen, sätter du textmarkören i dokumentet och använder Ångra-funktionen (via Redigera -menyn eller tangentbordet).  
Det går även att kopiera åt motsatt håll via dra-och-släpp:  
En texttabell eller ett markerat område i ett tabelldokument kan dras via dra-och-släpp till en tabellcontainer i Explorer för datakällor.  
Enkel text kan kopieras från ett dokument till ett datafält via dra-och-släpp.  
Anvisningar om detta finns i %PRODUCTNAME -hjälpen.  
Överföra data till ett textdokument  
Du kan infoga ett databasfält i ett textdokument genom att med musen dra ett fältnamn från kolumnhuvudet i datakällvyn till dokumentet.  
Då infogas ett fältkommando för det här databasfältet i dokumentet.  
Detta är mycket praktiskt när du skapar standardbrev (kopplad utskrift).  
Dra önskade fält för adress, tilltal o.s.v. till dokumentet.  
Det bästa sättet att infoga en komplett datapost är att markera motsvarande radhuvud och dra det till dokumentet.  
När du sedan släpper musknappen visas dialogrutan Infoga databaskolumner.  
Här kan du bestämma om alla databasfält ska tas med och om data ska kopieras till dokumentet i form av text, tabell eller fält.  
Alla dataposter som är markerade infogas.  
Överföra data till ett tabelldokument  
I ett tabelldokument kan du infoga en eller flera dataposter i den aktuella tabellen genom att markera raderna i datakällvyn och dra och släppa dem i tabelldokumentet.  
Data infogas på den plats där du släpper musknappen.  
Infoga kontrollfält i ett textformulär  
Om du utformar ett textformulär som är kopplat till en databas kan du skapa kontrollfält via dra-och-släpp från datakällvyn:  
Om du drar en databaskolumn till textdokumentet infogas ett fältkommando.  
Om du håller ner Skift + Kommando Ctrl när du drar infogas ett textfält grupperat med ett tillhörande etikettfält.  
Textfältet innehåller redan all databasinformation som du behöver till formuläret.  
Kopiera grafik från Gallery  
Dra ett grafikobjekt från Gallery till ett text-, tabell - eller presentationsdokument, så infogas grafikobjektet där.  
Om du släpper grafikobjektet direkt på ett ritobjekt gäller följande:  
Om objektet flyttas (dra utan att hålla ner någon tangent, inget särskilt tecken visas vid muspekaren) överförs bara teckenattributen från grafikobjektet och tilldelas ritobjektet som du släpper musknappen på.  
Om det kopieras (håll ner Ctrl-tangenten och dra, ett plustecken visas vid muspekaren) infogas grafikobjektet som objekt.  
Om en hyperlänk skapas (håll ner Skift+Ctrl-tangenterna och dra, en länkpil visas vid muspekaren) ersätts ritobjektet med grafikobjektet från Gallery, men det ersatta ritobjektets position och storlek bibehålls.  
Så här infogar du grafik från ett dokument till Gallery  
Du kan överföra ett intressant grafikobjekt, t.ex. från en HTML-sida, till Gallery genom att använda dra-och-släpp.  
Visa Gallery-temat där du vill placera grafikobjektet.  
Peka på grafikobjektet med musen utan att klicka.  
Om muspekaren förvandlas till en handsymbol är en hyperlänk kopplad till grafikobjektet.  
I så fall måste du hålla ner Alternativ Alt -tangenten när du klickar på grafikobjektet för att markera det utan att hyperlänken aktiveras.  
Om muspekaren inte förvandlas till en handsymbol, klickar du helt enkelt på grafikobjektet så att det markeras.  
Sedan klickar du på nytt på grafikobjektet och håller ner musknappen i minst två sekunder utan att flytta på musen.  
Då kopieras grafikobjektet till ett internminne.  
Dra nu grafikobjektet, utan att släppa musknappen, till Gallery.  
Ritobjekt som du har skapat med utrullningslisten Ritfunktioner kan inte läggas till i Gallery.  
Kopiera grafik mellan dokument  
Om du vill infoga ett grafikobjekt från ett dokument till ett annat dokument, kan du kopiera grafikobjektet genom att använda dra-och-släpp.  
Om du vill publicera ditt dokument bör du följa lagen om upphovsrätt och inhämta tillstånd från författarna till originalsidan för säkerhets skull.  
Öppna dokumentet där du vill infoga grafikobjektet.  
Öppna dokumentet som du vill kopiera grafikobjektet från.  
Håll ner Alternativ Alt -tangenten och klicka på grafikobjektet så att det markeras, men så att en hyperlänk som eventuellt är kopplad till det inte aktiveras.  
Håll ner musknappen och vänta ett ögonblick medan grafikobjektet kopieras till urklippet.  
Dra grafikobjektet till det andra dokumentet.  
Om dokumenten inte är synliga bredvid varandra, drar du först muspekaren till måldokumentets kommandoknapp.  
Fortsätt att hålla ner musknappen!  
Dokumentet aktiveras och visas och du kan föra muspekaren till dokumentet.  
Släpp musknappen så snart den gråa textmarkören antyder önskad plats för infogning av grafikobjektet.  
En kopia av grafikobjektet infogas.  
Om grafikobjektet är kopplat till en hyperlänk infogas hyperlänken i stället för grafikobjektet.  
Kopiera tabellområde till textdokument  
Öppna textdokumentet och tabelldokumentet.  
Markera det tabellområde som du vill kopiera.  
Peka i det markerade området, tryck på musknappen och håll ner den, vänta ett ögonblick och dra sedan området till textdokumentet.  
Om dokumenten inte är synliga bredvid varandra, drar du först muspekaren till måldokumentets kommandoknapp.  
Fortsätt att hålla ner musknappen!  
Dokumentet aktiveras och visas och du kan föra muspekaren till dokumentet.  
Släpp musknappen så snart textmarkören antyder platsen där du vill infoga tabellområdet.  
Tabellområdet infogas som OLE-objekt.  
Du kan när som helst markera och redigera OLE-objektet.  
Om du vill redigera OLE-objektet räcker det att dubbelklicka på det.  
Alternativt kan du markera objektet och välja Redigera - Objekt - Redigera eller Redigera på snabbmenyn.  
Objektet redigeras i en egen ram i textdokumentet, men du ser ikonerna och menykommandona som används för tabelldokument.  
Du öppnar OLE-objektets källdokument med kommandot Öppna.  
Dra-och-släpp inom %PRODUCTNAME -dokument  
Det finns många sätt att flytta eller kopiera objekt med dra-och-släpp.  
Markerad text, textområden, ritobjekt, grafik, kommandoknappar och andra formulärfunktioner, hyperlänkar, tabellområden och mycket annat går att flytta med musen.  
Var alltid uppmärksam på muspekaren när du drar.  
Den visar ett plustecken vid kopiering och en pil när en länk eller hyperlänk skapas.  
Muspekare  
Betydelse  
Flytta  
Kopiera  
Skapa en länk  
Om du håller ner Ctrl-tangenten eller Skift+Ctrl när du släpper musknappen, kan du oftast påverka om ett ojekt kopieras, flyttas eller om en länk skapas.  
Om du drar objekt från Navigator definierar du på undermenyn till ikonen Draläge om objektet kopieras eller om en länk eller en hyperlänk infogas.  
Om du har påbörjat en dra-och-släpp-aktivitet kan du avbryta den genom att trycka på Esc-tangenten innan du släpper musknappen.  
Ändra symbollist  
Om du t.ex. vill kopiera en ikon från en objektlist till funktionslisten, så att ikonen alltid är synlig, håller du bara ner Alt-tangenten och drar ikonen till sin nya plats. %PRODUCTNAME kommer automatiskt ihåg vad symbollisterna innehåller.  
Om du vill radera en ikon håller du ner Alt-tangenten och drar den från dess symbollist och släpper den utanför symbollisten.  
Om du vill ha ett streck på symbollisten drar du en ikon lite åt höger samtidigt som du håller ner Alt-tangenten.  
För att radera ett streck håller du ner Alt-tangenten och drar ikonen till höger om strecket lite åt vänster.  
På symbollisternas snabbmeny hittar du kommandot Synliga knappar.  
Med det öppnas en undermeny med en lista över de fördefinierade ikonerna.  
Ikoner som är markerade med en bock är synliga på symbollisten.  
Klicka på en post för att växla från synlig ikon till dold och tillbaka.  
Använd också kommandot Synliga knappar på en snabbmeny till en symbollist för att få en snabb översikt över namnen på ikonerna och deras funktioner.  
Skicka dokument som e-post  
Du kan skicka det aktuella dokumentet som bilaga till ett e-brev.  
Välj Arkiv - Skicka - Dokument som e-post.  
%PRODUCTNAME öppnar ditt standardprogram för e-post.  
Om du vill använda ett annat program, väljer du ut det under Verktyg - Alternativ - %PRODUCTNAME - Hjälpprogram.  
I ditt e-postprogram anger du en mottagare, ett ämne och skriver mer text om du vill och skickar iväg e-brevet.  
Hjälpprogram  
Spara dokument i externt format (t.ex. Microsoft)  
Välj kommandot Arkiv - Spara som.  
Dialogrutan Spara som öppnas.  
I fältet Filtyp väljer du ett externt format.  
Ange ett namn i fältet Filnamn och klicka på Spara.  
Om du alltid vill spara dina %PRODUCTNAME -dokument i ett externt format, väljer du det under Verktyg - Alternativ - Ladda / spara - Allmänt i området Standardfilformat.  
Spara som  
Sända fax och konfigurera %PRODUCTNAME för faxning  
Om du vill skicka ett fax direkt från %PRODUCTNAME behöver du ett faxmodem och en faxdrivrutin, som tillåter program att använda faxmodemet som en skrivare.  
Så här skickar du ett fax via en dialogruta  
Skriv ut det aktuella dokumentet med faxen som skrivare.  
Öppna dialogrutan Skriv ut genom att välja Arkiv - Skriv ut och välj faxdrivrutinen i kombinationsfältet Namn.  
När du klickar på OK öppnas en dialogruta för faxdrivrutinen där du kan ange faxmottagare.  
Så här konfigurerar du %PRODUCTNAME för faxning via en ikon  
Du kan konfigurera faxning från %PRODUCTNAME så att du bara behöver klicka på en ikon när du vill skicka iväg ett fax:  
Öppna Verktyg - Alternativ - Textdokument - Skriv ut.  
Välj faxdrivrutin i kombinationsfältet Fax och stäng dialogrutan med OK.  
Öppna snabbmenyn på funktionslisten och klicka på Synliga knappar.  
Du ser en lista med ikoner som kan konfigureras direkt för den här symbollisten.  
Alla ikoner som visas är markerade.  
Markera ikonen Skicka standardfax på snabbmenyn genom att klicka på den.  
Ikonen är nu synlig på funktionslisten.  
Om du klickar på ikonen startas faxdrivrutinen som du angav i steg 2 så att du kan faxa det aktuella dokumentet.  
Ändra ikonvy  
Du kan växla mellan flata ikoner och 3D-ikoner.  
Välj Verktyg - Alternativ - %PRODUCTNAME.  
Klicka på Vy och ta bort markeringen framför Flata ikoner.  
Klicka på OK.  
Med rutan Flata ikoner kan du byta mellan flat vy och 3D-vy.  
Med rutan Stora ikoner byter du mellan stora och små ikoner.  
Använda utrullningslist  
På verktygslisten till ett textdokument ser du ikonen Infoga längst upp.  
Du ser att ett fönster öppnas som innehåller fler ikoner.  
Du kan nu välja att antingen klicka på ikonen som du vill aktivera, eller att placera musen på utrullningslistens titellist och dra bort den från verktygslisten med nertryckt musknapp (du måste släppa musknappen en gång innan, annars kan du inte placera musen på titellisten).  
Lägg märke till ikonen på verktygslisten med vilken du öppnade utrullningslisten.  
Där ser du alltid den ikon som du har använt senast.  
Om du t.ex. klickar på ikonen Infoga grafik visas den här ikonen även på verktygslisten.  
Om du klickar kort på ikonen aktiverar du den funktion som är direkt synlig, om du klickar längre öppnas utrullningslisten igen.  
Symbollister vid textdokument  
Infoga och redigera kommandoknapp  
Öppna utrullningslisten Formulärfunktioner.  
Klicka på ikonen Kommandoknapp i utrullningslisten Formulär.  
Markören blir nu till ett hårkors.  
Kvadraten anger var kommandoknappen ska placeras och hur stor den ska vara.  
Den nya kommandoknappen är markerad.  
Du kan också hålla ner Alternativ Alt -tangenten samtidigt som du klickar.  
En markerad kommandoknapp kan du flytta och ändra storlek på precis som ett grafikobjekt.  
Via kommandoknappens snabbmeny kan du öppna dialogrutor där du redigerar kommandoknappens egenskaper.  
Välj Kontrollfält på snabbmenyn till den markerade kommandoknappen.  
Kommandoknapp visas.  
Du kan också öppna dialogrutan genom att klicka på knappen Kontrollfältegenskaper på utrullningslisten Formulärfunktioner.  
I den här dialogrutan kan du ändra texten på kommandoknappen under Allmänt - Rubrik.  
Om du vill att ett makro skall köras när du klickar på kommandoknappen anger du detta under fliken Händelser.  
När du klickar på någon av kommandoknapparna med tre punkter öppnas dialogrutan Tilldela makro.  
I listrutan Händelse listas samtliga händelser som kan kopplas till kommandoknapparna.  
Välj ett makro som skall köras när du klickar på kommandoknappen.  
Klicka sedan på Tilldela.  
Avsluta utkastläget med ikonen på utrullningslisten Formulärfunktioner.  
Om du nu klickar på kommandoknappen (inte på kanten) i dokumentet körs det tilldelade makrot.  
Förutom det markerade kontrollfältets egenskaper kan du också kontrollera egenskaperna hos det formulär som kontrollfältet tillhör.  
Klicka på ikonen Formuläregenskaper på utrullningslisten Formulär.  
I formuläret definieras bl.a. med vilken databas och tabell som kontrollfälten i formuläret ska kopplas ihop.  
Även för formuläret kan du koppla samman händelser med makron.  
Välj fliken Händelser.  
Här kan t.ex. alltid ett visst makro aktiveras när formuläret laddas.  
De övriga symbolerna på utrullningslisten Formulärfunktioner används till att definiera egna interaktiva dokument.  
I %PRODUCTNAME Basic kan du dessutom definiera egna dialogrutor - till detta finns det några fler kontrollfält för dialogrutor i %PRODUCTNAME Basic-IDE.  
Infoga, flytta och radera ikon på symbollist  
Beskrivningen gäller för alla funktioner som är möjliga i %PRODUCTNAME (inklusive egna makron).  
Öppna ett dokument av den typ som du vill ändra symbollisten för.  
Om du t.ex. vill ändra textobjektlisten för alla textdokument öppnar du ett textdokument.  
Öppna symbollistens snabbmeny och välj Redigera.  
Välj kategori och funktion i den nedre delen av dialogrutan.  
Om du inte hittar någon passande ikon för den här funktionen klickar du på Ikoner... och väljer en ikon.  
Bekräfta med OK.  
Dra nu den valda ikonen med nertryckt musknapp från dialogrutan till symbollisten.  
Släpp musknappen där du vill placera den nya ikonen.  
Stäng dialogrutan.  
Om du vill flytta den här ikonen till en annan plats, håller du ner Alternativknappen Alt-tangenten och drar ikonen dit du vill ha den (bara möjligt i Windows).  
Om du vill ta bort en ikon från symbollisten håller du ner Alternativknappen Alt-tangenten och drar bort ikonen från symbollisten (bara möjligt i Windows).  
Om symbollisten ska förankras vid en annan kant gör du så här:  
Håll ner Ctrl-tangenten och dubbelklicka på ett grått område på symbollisten.  
Den blir ett fritt fönster.  
Dra symbollisten till dess nya plats.  
Om du håller ner Ctrl-tangenten när du släpper musknappen och symbollisten är placerad ovanför en fönsterkant förankras symbollisten vid fönsterkanten.  
Verktyg - Anpassa  
Infoga ett objekt från Gallery  
Du kan antingen infoga ett objekt som Kopia eller som Länk i ett dokument.  
Kopian av ett objekt är oberoende av det ursprungliga objektet.  
Ändringar av originalobjektet påverkar inte kopian.  
Ändringar av originalobjektet påverkar även länken.  
Infoga ett objekt som kopia  
Öppna Gallery.  
Välj ett tema i det vänstra området.  
Markera objektet genom att klicka på det.  
Dra objektet till dokumentet eller öppna snabbmenyn genom att klicka med höger musknapp och välj Lägg till och Kopia.  
Infoga ett objekt som länk  
Öppna Gallery.  
Välj ett tema i det vänstra området.  
Markera objektet genom att klicka på det.  
Håll ner Skift+Ctrl-tangenterna och dra objektet till dokumentet eller öppna snabbmenyn genom att klicka med höger musknapp och välj Lägg till och Länk.  
Infoga ett objekt som bakgrundsgrafik  
Öppna Gallery.  
Välj ett tema i det vänstra området.  
Markera objektet genom att klicka på det.  
Öppna snabbmenyn och välj Lägg till - Bakgrund - Sida eller Stycke.  
Infoga ett objekt som textur (mönster) för ett andra objekt  
Öppna Gallery.  
Välj ett tema i det vänstra området.  
Markera objektet genom att klicka på det.  
Håll ner Ctrl-tangenten och dra objektet till det andra objektet i dokumentet.  
Redigera hyperlänk  
Så här ändrar du hyperlänktexten  
Möjlighet 1: håll ner Alternativ Alt -tangenten och klicka på hyperlänken.  
Möjlighet 2: klicka på fältet HYP på statuslisten så att SEL står där.  
Möjlighet 3: flytta markören till hyperlänken med piltangenterna.  
Nu kan du redigera texten utan att hyperlänken utförs.  
Så här ändrar du en hyperlänks URL  
Möjlighet 1: flytta markören till hyperlänken och öppna Hyperlnk-dialogrutan (ikon på funktionslisten).  
Möjlighet 2: öppna Hyperlänklisten (Visa - Symbollister - Hyperlänklist).  
Klicka på hyperlänken, släpp inte musknappen och dra hyperlänken till hyperlänklisten.  
Muspekaren visar var du kan släppa hyperlänken.  
Redigera URL:en på hyperlänklisten och tryck på Retur.  
Så här ändrar du attributen för alla hyperlänkar  
Du redigerar färg och formatering för hyperlänkar i ditt dokument via teckenformatmallarna "Internetlänk" och "Använd Internetlänk "i Stylist.  
Så här redigerar du en hyperlänk i form av kommandoknapp  
Om hyperlänken har formen av en kommandoknapp, så klickar du på kanten, eller så håller du ner Alternativ Alt -tangenten när du klickar på kommandoknappen.  
Den markeras då, och du kan öppna dialogrutan Egenskaper: Kommandoknapp  
Där kan du redigera den synliga texten under "Etikett" och URL:en under "URL ".  
Så här stänger du av den automatiska igenkänningen av hyperlänkar  
De automatiska igenkänningen av hyperlänkar stänger du av och sätter på under Verktyg - AutoKorrigering / AutoFormat - Alternativ i rutan Känn igen URL.  
Infoga hyperlänk  
Du kan infoga hyperlänkarna på två sätt: som text eller som kommandoknapp.  
I båda fallen kan den synliga texten skilja sig från URL:en.  
Du öppnar hyperlänklisten genom att välja Visa - Symbollister - Hyperlänklist.  
I det vänstra fältet matar du in den synliga texten, i det högra fältet den fullständiga URL:en, inklusive http: / / eller file: / /.  
Placera textmarkören på det ställe där hyperlänken ska infogas i dokumentet.  
Klicka sedan på ikonen Länk på hyperlänklisten resp. på Överta i hyperlänkdialogrutan.  
Hyperlänken infogas som text.  
Om du vill infoga hyperlänken som kommandoknapp, håller du ner musknappen något längre på ikonen Länk, och väljer Som knapp på undermenyn resp. väljer posten Knapp i fältet Form i hyperlänkdialogrutan.  
Om du i stället för hyperlänklisten hellre vill använda hyperlänk-dialogrutan för att definiera hyperlänken, kan du öppna den med ikonen på funktionslisten.  
Om du vill hoppa till ett visst ställe i samma textdokument, infogar du ett bokmärke på det stället (Infoga - Bokmärke).  
Om du vill göra en länk till en cell i en tabell, ger du cellen ett namn (Infoga - Namn - Definiera).  
I kombinationsfältet Samlingsbox till webbadresser matar du vid hopp inom samma dokument bara in URL:ens förkortning:  
Om bokmärket heter Hoppmål, matar du in #Hoppmål.  
Om du hoppar till ett annat dokument, matar du in den kompletta URL:en.  
Om du inte är så van vid URL-skrivsättet, kan du automatiskt få hjälp av %PRODUCTNAME: inmatningen C:\Doku\Fil1.sdw#Hoppmål ändrar %PRODUCTNAME automatiskt till det korrekt skrivna file: / //c _BAR_ / Doku / Fil1.sdw#Hoppmål.  
Hyperlänkar kan du även infoga genom att dra och släppa dem från Navigator.  
Hyperlänkarna kan hänvisa till referenser, överskrifter, grafik, tabeller, objekt, förteckningar eller bokmärken.  
Om du vill infoga en hyperlänk som hänvisar till Tabell 1 drar du posten Tabell 1 från Navigator till texten.  
Du måste ha valt draläget Infoga som hyperlänk i Navigator.  
Relativa och absoluta länkar  
Om du integrerar hyperlänkar, måste du ta hänsyn till (minst) två villkor, nämligen inställningen relativ / absolut när du sparar och frågan om filen finns eller inte:  
%PRODUCTNAME fungerar olika beroende på inställningen under Verktyg - Alternativ - Ladda / spara - Allmänt där du kan välja om länkarna ska skapas relativt eller absolut när de sparas.  
Relativ adressering är bara möjlig om utgångsdokumentet och målet för länken ligger på samma enhet.  
Du bör skapa samma katalogstruktur på din hårddisk som i ditt hemsida-område hos Internetleverantören.  
Kalla baskatalogen för din hemsida på din hårddisk för t.ex. "hemsida".  
Startfilen är då t.ex. "index.htm" med den kompletta sökvägsangivelsen "C:\homepage\index.htm ".  
På din leverantörs server kan det t.ex. bli följande URL: "http: / /www.minprovider.com / minsida / index.htm".  
Vid relativ adressering anger du länken relativt till utgångsdokumentets plats.  
Om du t.ex. har arkiverat all grafik på din hemsida i en underordnad mapp "C:\homepage\grafik", så anger du följande sökväg som mål för grafiken "bild.gif": "grafik\bild.gif".  
Det är den relativa sökvägen som utgår från platsen för filen "index.htm".  
På leverantörens server lägger du bilden i mappen "minsida / grafik". %PRODUCTNAME kommer automatiskt att kopiera grafiken till rätt katalog på servern om du överför dokumentet "index.htm" via dialogrutan Arkiv - Spara som till leverantörens server, och om du har markerat rutan Kopiera lokal grafik till Internet under Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet.  
En absolut sökväg som "C:\homepage\grafik\bild.gif" skulle inte längre fungera på leverantörens server.  
Varken på servern eller på datorn hos en läsare av din Internetsida måste det finnas en enhet C: (operativsystem som Unix eller MacOS har inga enhetsbokstäver), och även om mappen homepage\grafik fanns där, så skulle inte Din bild finnas där.  
Använd alltså hellre relativ adressering för fillänkar.  
En länk på en annan webbsida som t.ex. "www.sun.se" eller "www.minleverantör.com / minsida / index.htm "är en absolut länk.  
%PRODUCTNAME fungerar också olika beroende på om filen som länken refererar till finns eller inte finns och var den finns. %PRODUCTNAME kontrollerar varje ny länk och sätter automatiskt in mål och protokoll.  
Resultatet ser du i den skapade HTML-koden när du har sparat utgångsdokumentet (inte i länkens tipshjälp, se nedan).  
Följande regler gäller:  
En relativ adressering ("grafik / bild.gif") är bara möjlig om båda filerna finns på samma enhet.  
Om båda filerna finns på olika enheter, men i lokala filsystem, sker en absolut adressering med "file :"-protokoll ("file: / //data1 / xyz / bild.gif").  
Om båda filerna finns på olika servrar eller om målet för länken inte finns för närvarande, sker en absolut adressering med "http :"-protokoll ("http: / /data2 / abc / bild.gif").  
Se alltså till att du ordnar alla filer som du behöver på din hemsida på samma enhet som hemsidans startfil.  
På det här sättet kan %PRODUCTNAME automatiskt sätta in protokollet och målet så att referensen även fungerar på leverantörens server.  
I tipshjälpen till en hyperlänk och i HTML-källtextsredigeraren ser du alltid det absoluta skrivsättet eftersom %PRODUCTNAME alltid arbetar med absoluta sökvägar internt.  
Vad som skrivs i filen vid HTML-export ser du först när du tittar på resultatet av HTML-exporten, t.ex. genom att du laddar den skapade HTML-filen som "Text" eller öppnar den med en texteditor.  
Söka med hyperlänklisten  
Sökning med hyperlänklisten beskrivs utförligt i %PRODUCTNAME -hjälpen.  
Skriv den text som du söker efter i fältet URL-namn.  
Om du dubbelklickar på ett ord i texten förs det in automatiskt.  
Öppna undermenyn till ikonen Sök genom att klicka på den.  
Välj den önskade sökmotorn genom att klicka på den.  
%PRODUCTNAME öppnar din webbläsare och den upprättar förbindelsen till sökmotorn.  
Efter en stund visas sökresultatet på bildskärmen.  
Hyperlänklist  
Öppna dokument i externt format (t.ex. Microsoft)  
Öppna ett dokument i ett externt format då och då  
Välj Arkiv - Öppna.  
I fältet Filtyp väljer du ett externt format.  
Välj ett namna och klicka på Öppna.  
Öppna dokument i ett externt format ofta  
Om du alltid vill öppna dina dokument i ett externt format, väljer du det under Verktyg - Alternativ - Ladda / spara - Allmänt i området Standardfilformat.  
Konvertera alla dokument i en mapp  
Öppna AutoPiloten som hjälper dig att konvertera alla dokument från Microsoft Word, Microsoft Excel eller Microsoft Powerpoint till %PRODUCTNAME -dokument.  
Du kan välja käll - och målkatalog, om du vill konvertera dokument och / eller dokumentmallar, med mera.  
Välj Arkiv - AutoPilot - Dokumentkonverterare.  
Arbeta med VBA-kod  
Infoga, redigera och spara bitmap  
Infoga bitmap  
En bitmapbild kan infogas i dokument från %PRODUCTNAME Writer, %PRODUCTNAME Calc, %PRODUCTNAME Draw och %PRODUCTNAME Impress.  
Välj Infoga - Grafik - Från fil.  
I %PRODUCTNAME Draw och %PRODUCTNAME Impress heter kommandot Infoga - Grafik.  
Välj ut en fil.  
Med fältet Filtyp kan du begränsa urvalet till vissa filtyper.  
Markera rutan Länka om du vill ha en länk till originalfilen.  
Om rutan Länka är markerad laddas bitmapbilden om varje gång du uppdaterar och laddar dokumentet, sedan används redigeringsstegen som du har gjort på den lokala kopian av bilden igen och bilden visas.  
Om rutan Länka inte är markerad, arbetar du alltid bara med kopian som skapades när bilden infogades i dokumentet första gången.  
Klicka på Öppna för att infoga bilden.  
Redigera bitmap  
Om du markerar bitmapbilden innehåller objektlisten verktygen som du behöver om du vill redigera bilden.  
Det är alltid bara en lokal kopia som redigeras i dokumentet, även om du har infogat en bild som länk.  
Objektlistens utseende kan variera något beroende på med vilken modul du arbetar.  
Illustrationen visar objektlisten i %PRODUCTNAME Draw objektlisten i %PRODUCTNAME Draw objektlisten i %PRODUCTNAME Draw:  
Det finns ett antal filter på utrullningslisten Filter som du öppnar med ikonen längst till vänster på objektlisten:  
När du klickar på några av filtren öppnas en dialogruta där du t.ex. kan välja intensitet för filtret.  
Du kan förse bitmapbilden med text och grafik, markera de här objekten tillsammans och exportera markeringen som en ny bitmapbild.  
Spara bitmap  
Om du vill spara ändringarna av en bitmapbild som bildfil, t.ex. i filformatet GIF, JPEG eller TIFF, måste du markera och exportera bitmapbilden.  
Detta kan du bara göra i %PRODUCTNAME Draw och %PRODUCTNAME Impress.  
Markera bitmapbilden.  
Markera eventuellt även andra objekt (håll ner skifttangenten när du markerar eller rita upp en ram runt alla objekt) om du t.ex. vill förse bitmapbilden med text.  
Välj Arkiv - Exportera.  
Dialogrutan Exportera visas.  
Välj filformat i fältet Filtyp, t.ex. GIF eller JPEG.  
Om du bara vill exportera de markerade objekten, markerar du rutan Markering.  
Om Markering inte är markerad exporteras hela dokumentsidan.  
Ange ett namn för filen och klicka på Spara.  
Rita ett grafikobjekt med ritfunktionerna  
Öppna Ritfunktionerna på verktygslisten.  
Om du har valt en funktion visas motsvarande ikon på verktygslisten.  
Om du klickar längre öppnas utrullningslisten där du kan välja en annan funktion.  
Ritobjekt går att redigera och ändra i efterhand.  
Vid sådana teckningselement rör det sig om vektorgrafik som du kan skala som du vill utan kvalitetsförlust.  
Dra utrullningslisten som eget fönster till bildskärmen om du vill rita flera element.  
Du skapar en rektangel genom att klicka på rektangelikonen och sedan peka på den plats i dokumentet där ett hörn av rektangeln ska placeras.  
Tryck på musknappen här, håll ner den och dra till motstående hörnet av rektangeln.  
Om du släpper musknappen infogas rektangeln i dokumentet.  
Den är markerad och du kan redigera dess egenskaper via snabbemenyn.  
Om du inte vill rita upp ritobjektet från ett hörn till det motstående hörnet utan från mitten, håller du ner Alternativ Alt -tangenten.  
Om du håller ner skifttangenten när du drar begränsar du det skapade objektet, i stället för en rektangel med olika långa sidor ritas t.ex. en kvadrat upp.  
Om du vill skala objekten markerar du dem först genom att klicka på dem med urvalsverktyget.  
Då ser du åtta handtag runt objektet.  
Om du drar ett av de fyra handtagen i hörnen fixeras det motstående hörnet, medan det går att flytta de andra tre hörnen.  
Om du drar ett av de fyra handtagen mitt på sidorna, fixeras den motstående sidan.  
Om du vill flytta ritobjekt markerar du dem först (en och en eller flera samtidigt genom att hålla ner skifttangenten).  
Textobjekt markerar du genom att klicka på deras kant.  
Sedan håller du ner musknappen och drar objekten till den nya platsen.  
Om du håller ner skifttangenten när du drar så kan du bara placera objekten på vissa ställen som är orienterade efter sidmarginalerna och de andra objekten på sidan.  
Om du håller ner Kommando Ctrl -tangenten när du drar ritobjektet kopieras det.  
När du har skapat och redigerat ritobjekt återvänder du till det normala textläget genom att klicka på ett området i dokumentet där inga ritobjekt eller andra objekt finns.  
Om du är i ett ritläge avslutar du det först genom att t.ex. klicka på ikonen Urval.  
Information om de olika ikonerna  
Infoga specialtecken  
Så här infogar du specialtecken (t.ex. bockar, rutor, telefonsymboler) i din text.  
Välj Infoga - Specialtecken så att du kan välja bland alla tecken.  
Klicka på ett eller flera tecken efter varandra i det stora urvalsfältet.  
Tecknen visas vid den undre kanten av dialogrutan.  
Stäng dialogrutan med OK så infogas alla visade tecken med det valda teckensnittet i det aktuella dokumentet.  
Dialogrutan Specialtecken kan du öppna i alla textinmatningsfält (t.ex. i URL-fältet på funktionslisten, i inmatningsfälten i Sök och ersätt-dialogrutan o.s.v.) genom att trycka Skift + Kommando Ctrl +S.  
Det finns för närvarande bara tre möjligheter att mata in bokstäver med accent direkt från tangentbordet.  
Sun Solaris: använd ett Sun-tangentbord.  
Tryck först på Compose-tangenten till höger om blanksteg, sedan matar du in den första och andra modifiern.  
Linux / NetBSD: använd dead-keys.  
Tryck först på tangenten ´ eller ` i ett xterm-fönster.  
Tecknet får inte synas på bildskärmen.  
Tryck nu t.ex. på e.  
E:et får en accent som é eller è.  
Ersätt i så fall den.  
Eventuellt kan du också ha satt miljövariabeln SAL_NO_DEADKEYS som stänger av dead-keys.  
AltGr som extra Compose-tangent.  
Tangenten AltGr kan arbeta som Compose-tangenten i %PRODUCTNAME om du sätter miljövariabeln SAL_ALTGR_COMPOSE.  
AltGr-tangenten måste utlösa en Mode_switch, alltså måste t.ex. xmodmap -e "keysym Alt_R = Mode_switch" vara satt.  
Tryck först på AltGr, sedan den första modifiern, sedan den andra modifiern.  
Tecknen sammanfogas så som är beskrivet i filen / usr / openwin / include / X11 / Suncompose.h i ett Solarissystem.  
Specialtecken  
Ändra en installation  
Du kan anpassa en installation av %PRODUCTNAME i efterhand genom att lägga till nya och ta bort installerade komponenter.  
Starta Setupprogrammet för %PRODUCTNAME antingen via Windows-startmenyn eller antingen via startlisten eller direkt från installationskatalogen för %PRODUCTNAME.  
{installdir}\program\setup.exe {installdir} / setup  
{installdir} betecknar katalogen där du har installerat %PRODUCTNAME.  
Välj Modifiera som installationsalternativ från installationsdialogrutan och följ anvisningarna på bildskärmen.  
I de följande dialogrutorna kan du välja ut vilka komponenter som ska installeras eller avinstalleras.  
Reparera en skadad installation  
Om delar av %PRODUCTNAME inte längre fungerar som de ska på grund av skadade programfiler eller registreringsposter, kan du reparera installationen med hjälp av setupprogrammet.  
Starta Setupprogrammet för %PRODUCTNAME antingen via Winows-startmenyn eller antingen via startlisten eller direkt från installationskatalogen för %PRODUCTNAME.  
{installpath}\program\setup.exe {installpath} / setup  
{installdir} betecknar katalogen där du har installerat %PRODUCTNAME.  
Välj Reparera som installationsalternativ från installationsdialogrutan och följ anvisningarna på bildskärmen.  
Skriva ut etiketter med adresser  
Om du vill skapa adressetiketter, t.ex. för standardbrev (kopplad utskrift) som inte passar i fönsterkuvert, gör du så här:  
1.  
Öppna via Arkiv - Nytt - Etiketter dialogrutan Etiketter.  
2.  
Välj formatet för etikettarken som du vill skriva ut.  
Tänk på att rutan Synkronisera innehåll måste vara förkryssad under fliken Tillägg.  
Stäng dialogrutan med Nytt dokument.  
3.  
När du ser etikettdokumentet öppnar du datakällvyn genom att trycka på F4.  
Klicka på nålsymbolen i kanten av datakällvyn om den täcker den första etiketten.  
4.  
Välj tabellen från din adressdatakälla i datakällvyn.  
5.  
Dra datafälten som behövs i adressen en och en till etiketten uppe till vänster.  
Klicka t.ex. på kolumnhuvudet NAME, håll ner musknappen och dra till etiketten.  
Ett fältkommando infogas.  
Placera fältkommandona för den fullständiga adressen på den första etiketten uppe till vänster.  
6.  
Sätt markören vid den sista textpositionen (efter det sista fältkommandot) på den första etiketten.  
7.  
Öppna dialogrutan Fältkommandon, t.ex. med tangentkombinationen Kommando Ctrl +F2, och klicka på fliken Databas.  
8.  
Välj fälttypen Nästa datapost, klicka på Infoga och Stäng.  
9.  
Nu kan du synkronisera etiketterna.  
Klicka på kommandoknappen Synkronisera i det lilla fönstret.  
10.  
I datakällvyn markerar du dataposterna som du vill ha på adressetiketterna genom att klicka på radhuvudena.  
Använd Skift - eller Kommando Ctrl -tangenten på det vanliga sättet för att markera flera dataposter tillsammans.  
11.  
Klicka på ikonen Data i fält på Databaslisten.  
12.  
Sedan kan du spara och / eller skriva ut etikettdokumentet.  
Efter den sista etiketten på en sida utförs kommandot Nästa datapost automatiskt!  
Infoga alltså inte det här kommandot manuellt efter den sista etiketten på en sida.  
Skriva ut etiketter med löpande nummer  
Om du t.ex vill skriva ut lotter eller inträdesbiljetter med löpande nummer, gör du så här:  
Välj Arkiv - Nytt - Etiketter.  
Dialogrutan Etiketter öppnas.  
Välj ett format som du vill skriva ut under fliken Etiketter i området Format.  
De färdiga etikettarken eller rullarna som finns att köpa består oftast av starkare papper som är perforerat, eller av självhäftande lappar.  
Om du vill bestämma formatet själv kan du göra detta under fliken Format.  
Markera rutan Synkronisera innehåll under fliken Tillägg.  
Klicka på Nytt dokument.  
Det skapas nu ett nytt dokument med uppdelningen som du har valt.  
Du behöver bara redigera etiketten uppe till vänster och sedan trycka på kommandoknappen Synkronisera etiketter så att alla etiketter ser likadana ut.  
Kommandoknappen är bara synlig om du har kryssat för rutan Synkronisera innehåll under fliken Tillägg.  
Mata in text på etiketten uppe till vänster och formatera teckensnittet som du vill.  
Du får ett löpande nummer genom att infoga ett fältkommando.  
Sätt markören på det ställe där numret ska visas.  
Tryck på Kommando Ctrl +F2 eller välj Infoga - Fältkommando - Andra.  
I dialogrutan Fältkommandon klickar du på fliken Variabler.  
Välj fälttypen Sätt variabel om den inte redan är markerad.  
Mata in ett valfritt namn för räknevariabeln i fältet Namn, t.ex. Nummer.  
För att variabeln skall höjas med 1 för varje etikett, matar du in följande formel i textfältet Värde:  
Nummer+1.  
Klicka på Infoga och stäng dialogrutan Fältkommandon.  
Klicka på Synkronisera etiketter.  
Nu kan du spara och skriva ut det färdiga dokumentet.  
Skapa och skriva ut etiketter och visitkort  
Utforma visitkort via dialogruta  
Om du väljer Arkiv - Nytt - Visitkort öppnas en dialogruta med flera flikar där du kan välja hur dina visitkort ska se ut.  
Utforma etiketter och visitkort  
Det finns ett annat sätt att utforma visitkort: om man ser visitkort som ett specialfall av etiketter.  
Visitkort är i allmänhet likadana.  
Etiketter kan ha olika innehåll från en databas eller löpnummer.  
Välj Arkiv - Nytt - Etiketter, dialogrutan Etiketter öppnas.  
Klicka på fliken Etiketter och definiera etikettformatet i området Format.  
%PRODUCTNAME Writer innehåller många format från ark som finns att köpa färdiga med etiketter, visitkort och så vidare.  
Du kan lägga till användardefinierade format.  
Under fliken Etiketter väljer du etiketternas påskrift i området Påskrift.  
Det är ofta databasfält så att du kan skriva ut etikettsidorna med skiftande innehåll som "Standardbrev" (kopplad utskrift), men du kan också skriva ut samma text på alla etiketter.  
I kombinationsfälten väljer du ut databasen och tabellen som datafälten hämtas ifrån.  
Med pilknappen överför du det valda datafältet till påskriftsområdet.  
Du kan infoga en radbrytning med returtangenten och dessutom kan du mata in mellanslag och andra valfria fasta texter.  
Under fliken Format kan du definiera egna etikettformat som inte finns med bland de förinställda formaten.  
Förutsättningen för detta är att du har ställt in etikettypen "Användare" under fliken Etiketter.  
Under fliken Tillägg bestämmer du om alla etiketter eller bara vissa etiketter ska skapas.  
Rutan Synkronisera innehåll under fliken Tillägg är viktig.  
Om du markerar den behöver du bara mata in och redigera en etikett som ständigt återkommer en gång (i etiketten uppe till vänster).  
När du klickar på Nytt dokument öppnas ett litet fönster med kommandoknappen Synkronisera etiketter.  
Mata in den första etiketten.  
När du klickar på kommandoknapppen kopieras den aktuella enskilda etiketten till alla andra etiketter på arket.  
Klicka på Nytt dokument för att skapa ett nytt dokument med inställningarna som du har gjort.  
Skriv ut det nya dokumentet.  
Visitkort  
Välja språk i dokument  
Språket som du väljer för ditt dokument bestämmer bland annat vilken ordlista som används för rättstavningskontroll, synonymordlista och avstavning, vilka decimaltecken och tusentalsavgränsare som används och vilket valutaformat som är förinställt.  
I princip gäller språket som är inställt för hela dokumentet.  
Men inom dokumentet kan du tilldela varje styckeformatmall ett eget språk.  
Det har högre prioritet än språket för hela dokumentet.  
Inom ett stycke kan du tilldela utvalda textdelar ett språk, antingen som direkt formatering eller via en teckenformatmall.  
Den här tilldelningen har högre prioritet än styckeformatmall och dokumentspråk.  
Välja språk för hela dokumentet  
Välj Verktyg - Alternativ - Språkinställningar - Språk.  
I området Standardspråk för dokument väljer du dokumentspråk för alla nya dokument som du skapar.  
Om du markerar rutan Bara för det aktuella dokumentet gäller inställningen bara för det aktuella dokumentet.  
Stäng dialogrutan med OK.  
Välja språk för en styckeformatmall  
Placera markören i stycket vars styckeformatmall du vill redigera.  
Öppna snabbmenyn och välj Redigera styckeformatmall.  
Dialogrutan Styckeformatmall öppnas.  
Klicka på fliken Teckensnitt.  
Välj Språk och klicka på OK.  
Nu har alla stycken, som är formaterade med den aktuella styckeformatmallen, det valda språket.  
Tilldela markerad text språk direkt  
Markera texten som du vill tilldela ett språk.  
Välj Format - Tecken.  
Dialogrutan Tecken öppnas.  
Klicka på fliken Teckensnitt.  
Välj Språk och klicka på OK.  
I %PRODUCTNAME Calc väljer du Format - Cell och gör på samma sätt.  
Välja språk för teckenformatmall  
Öppna Stylist och klicka på ikonen Teckenformatmallar.  
Klicka på namnet på teckenformatmallen som ska få ett annat språk.  
Öppna snabbmenyn i Stylist och välj Ändra.  
Dialogrutan Teckenformatmall öppnas.  
Klicka på fliken Teckensnitt.  
Välj Språk och klicka på OK.  
Nu kan du tilldela den markerade texten teckenformatmallen.  
Verktyg - Alternativ - Språkinställningar - Språk  
Format - Tecken - Teckensnitt  
Allmänna anvisningar för %PRODUCTNAME  
Öppna och spara dokument och dokumentmallar  
Använda fönster, menyer, ikoner  
Kopiera data, med dra-och-släpp och per meny  
Datakällor  
Registrera ändringar (revideringsfunktion)  
Anpassa och ändra %PRODUCTNAME  
Diagram (charts)  
Övrigt  
Välja måttenheter  
Du kan välja måttenhet separat för %PRODUCTNAME Writer-, %PRODUCTNAME Writer / Web-, %PRODUCTNAME Calc-, %PRODUCTNAME Impress - och %PRODUCTNAME Draw-dokument.  
Välj Verktyg - Alternativ.  
Klicka på dokumenttypen som du vill välja måttenhet för.  
Klicka på Textdokument om du vill välja måttenhet för %PRODUCTNAME Writer.  
Klicka på Allmänt.  
Under Allmänt i området Inställningar finns det ett kombinationsfält där du kan välja måttenhet.  
Stäng dialogrutan med OK.  
Omräkning av måttenheter  
Verktyg - Alternativ - Textdokument - Allmänt  
Navigation för att snabbt komma till ett objekt  
Detta är den enklaste användningen av Navigator.  
Om du dubbelklickar på objektet i Navigator flyttas markören till objektens position i dokumentet.  
Du kan använda utrullningslisten Navigation till att bläddra till föregående eller nästa objekt i en viss kategori.  
Du öppnar utrullningslisten med ikonen Navigation nere till höger i dokumentfönstret eller uppe till vänster i Navigator.  
På utrullningslisten Navigation väljer du först kategori, sedan klickar du på en av ikonerna till höger, Föregående objekt eller Nästa objekt.  
Namnen på ikonerna rättar sig efter kategorin, ikonen för att bläddra vidare heter t.ex. beroende på kategori "Nästa sida" eller "Nästa bokmärke ".  
Navigator för överblick över dokumentet  
I det följande kallar vi för enkelhetens skull hela innehållet i Navigator-fönstret helt enkelt för "Kategori", oavsett om det är överskrifter, tabeller, textramar, grafiker, OLE-objekt, textramar, områden, hyperlänkar, referenser, mappar eller anteckningar.  
Navigator visar dig vilka kategorier som finns i dokumentet.  
Så snart du ser ett plustecken till vänster om namnet på kategorin, finns det minst ett objekt av detta slag.  
Hur många exakt ser du i den Aktiva hjälpen om du låter muspekaren stå kvar lite längre på namnet.  
Du öppnar en kategori genom att klicka på plustecknet.  
Om du bara är intresserad av posterna i den här kategorin kan du markera kategorin och klicka på ikonen Växla innehållsvisning.  
Då ser du bara objekten i den här kategorin tills du klickar på ikonen igen.  
Om fönstret i den förankrade Navigator är för litet kan du göra det till ett fritt fönster (håll ner Kommando Ctrl -tangenten och dubbelklicka på det gråa området).  
Då kan du ändra storleken hur du vill.  
Visa hjälpens navigationsområde  
I hjälpfönstret kan du visa eller dölja navigationsområdet efter behov:  
Klicka på ikonen till vänster på symbollisten i hjälpfönstret för att visa och dölja navigationsområdet.  
Så här stänger du av numrering / punktuppställning för enskilda stycken  
Om markören står i en numrering eller punktuppställning stänger du av den automatiska numreringen eller punktuppställningen i det aktuella stycket eller i de markerade styckena genom att klicka på ikonen Numrering av på numreringsobjektlisten respektive Numrering på / av på textobjektlisten.  
Om markören står i en numrering eller punktuppställning stänger du av den automatiska numreringen eller punktuppställningen i det aktuella stycket eller de markerade styckena genom att klicka på ikonen Punktuppställning på / av på objektlisten.  
Gör så här om du vill undanta ett stycke i en punktuppställning / numrering från den automatiska numreringen via tangentbordet:  
Ställ markören i början av ett numrerat stycke och tryck på backstegstangenten.  
Numreringen fortsätter i efterföljande stycke.  
Om du trycker på Retur i ett tomt numrerat stycke avslutas den aktuella numreringen.  
Format - Punktuppställning / numrering  
Välja maximalt möjligt sidformat  
Alla skrivare kan inte skriva ut ända ut i kanten.  
Men hur långt ut i kanten får egentligen texten eller grafiken gå för att allt skall få plats på sidan?  
%PRODUCTNAME ger dig en halvautomatisk hjälp som gör det möjligt för dig att skriva så långt ut i kanten som din skrivare tillåter.  
Kontrollera att rätt skrivare är inställd under Arkiv - Skrivarinställning....  
Kontrollera att onlinelayouten inte är aktiverad (i menyn Visa).  
Växla till fliken Sida.  
I området Marginaler kan du nu ställa in det maximala resp. det minimala värdet för de fyra marginalerna vänster, höger, övre och nedre, genom att trycka på tangenterna PageUp respektive PageDown.  
I förhandsvisningen ser du det utskrivbara området i form av en streckad rektangel.  
Stäng dialogrutan genom att klicka på OK.  
Skriva ut i svartvitt  
Om du har en färgskrivare men bara vill skriva ut i svartvitt finns det följande möjligheter:  
Skriva ut text och grafik i svartvitt  
Välj Arkiv - Skriv ut.  
Dialogrutan Skriv ut öppnas.  
Klicka på Egenskaper.  
Egenskapsdialogrutan för din skrivare öppnas.  
Välj alternativet för att skriva ut i svartvitt.  
Det finns mer information i hjälpen eller handboken till din skrivare.  
Bekräfta dialogrutan och klicka på OK i dialogrutan Skriv ut.  
Det aktuella dokumentet skrivs ut i svartvitt.  
Skriva ut i %PRODUCTNAME Impress och %PRODUCTNAME Draw  
Välj Verktyg - Alternativ - Presentation respektive Verktyg - Alternativ - Teckning.  
Klicka på Skriv ut.  
I området Utmatningskvalitet väljer du ett av alternativen Gråskalor eller Svartvitt och klickar på OK.  
Sedan skrivs alla presentationer respektive teckningar ut utan färg.  
Om du bara vill avstå från färg när du gör den aktuella utskriften, väljer du alternativet under Arkiv - Skriv ut - Fler.  
När du väljer alternativet Standard för utmatningskvaliteten skrivs färger ut igen.  
Gråskalor omvandlar allt till maximalt 256 steg från svart till vitt.  
Svartvitt omvandlar allt till de två värdena svart och vitt.  
Bara skriva ut text i svartvitt  
I %PRODUCTNAME Writer kan du välja att text som är formaterad i färg skrivs ut i svartvitt.  
Du kan välja mellan att definiera detta i förinställningarna för alla kommande textdokument som skrivs ut eller bara för en utskrift av det aktuella textdokumentet.  
Skriva ut alla textdokument med svartvit text  
Välj Verktyg - Alternativ - Textdokument eller Verktyg - Alternativ - HTML-dokument.  
Klicka på Skriv ut.  
Markera rutan Svart utskrift i området Innehåll och klicka på OK.  
Alla textdokument eller HTML-dokument skrivs nu ut med svart text.  
Skriva ut det aktuella textdokumentet med svartvit text  
Välj Arkiv - Skriv ut.  
Dialogrutan Skriv ut öppnas.  
Klicka på Fler.  
Dialogrutan Skrivaralternativ öppnas.  
Markera rutan Svart utskrift i området Innehåll och klicka på OK.  
Textdokumentet eller HTML-dokumentet som nu skrivs ut har svartvit text.  
Dialogrutan Skriv ut  
Dialogrutan Verktyg - Alternativ  
Skriva ut i annan ordningsföljd  
Så här skriver du ut dokument i rätt ordning.  
Välj Arkiv - Skriv ut och sedan kommandoknappen Fler.  
Bekräfta med OK.  
Nu skrivs den sista sidan ut först och den första sidan till sist.  
Skriv ut  
Skyddat innehåll i %PRODUCTNAME  
Här hittar du en översikt över de olika sätten att skydda innehåll i %PRODUCTNAME mot redigering, radering och visning.  
Skydda alla dokument som sparas  
Alla dokument som sparas i XML-format (%PRODUCTNAME 6.0-format), kan förses med ett lösenord.  
Utan lösenordet går det sedan inte att öppna dokumenten.  
Innehållet krypteras så att det inte heller går att läsa med en extern redigerare.  
Detta gäller för innehåll, grafik och OLE-objekt.  
Aktivera skydd  
Välj Arkiv - Spara som, markera rutan Spara med lösenord.  
Spara dokumentet.  
Avaktivera skydd  
Öppna dokumentet och mata in rätt lösenord.  
Välj Arkiv - Spara som, upphäv markering vid Spara med lösenord.  
Meta-informationen som du kan mata in under Arkiv - Egenskaper och som t.ex. innehåller ditt namn, skapandedatum, antal ord och tecken krypteras inte!  
Skydda revideringsfunktion  
Med revideringsfunktionen i %PRODUCTNAME Calc och %PRODUCTNAME Writer registreras vid varje ändring vem som har gjort ändringen.  
Den här funktionen kan aktiveras med skydd så att den bara går att stänga av om det riktiga lösenordet anges.  
Sålänge funktionen är aktiv registreras alla ändringar, att acceptera eller ignorera är inte möjligt.  
Aktivera skydd  
Välj Redigera - Ändringar - Skydda registrering.  
Ange ett lösenord som består av minst 5 tecken och bekräfta.  
Avaktivera skydd  
Välj Redigera - Ändringar - Skydda registrering.  
Ange rätt lösenord.  
Skydda cellområden i %PRODUCTNAME Calc  
I %PRODUCTNAME Calc kan du skydda hela tabeller och dokumentet i sin helhet.  
Då väljer du om cellerna ska skyddas mot oavsiktliga ändringar, om formlerna ska gå att se, om cellerna är synliga och / eller om cellerna ska kunna skrivas ut.  
Skyddet kan förses med ett lösenord men måste inte ha det.  
Om du har tilldelat ett lösenord kan skyddet bara upphävas när du har angett det korrekta lösenordet.  
Tänk på att cellskyddet för de celler som tilldelats attributet Skyddad först får effekt när du skyddar hela tabellen.  
I förinställningen har alla celler attributet Skyddad.  
Du upphäver alltså attributet för de celler där användaren får lov att göra ändringar.  
Sedan skyddar du hela tabellen och sparar dokumentet.  
Aktivera skydd  
För celler: markera cellområde.  
Välj Format - Cell - fliken Cellskydd.  
För tabeller: välj Verktyg - Skydda dokument - Tabell.  
För dokument: välj Verktyg - Skydda dokument - Dokument.  
Om du vill anger du ett lösenord som består av minst 5 tecken och bekräftar det.  
Avaktivera skydd  
För tabeller: välj Verktyg - Skydda dokument - Tabell.  
För dokument: välj Verktyg - Skydda dokument - Dokument.  
Om ett lösenord har tilldelats, ange rätt lösenord.  
Skydda textområden i %PRODUCTNAME Writer  
Alla områden i ett %PRODUCTNAME Writer-textdokument kan skyddas mot ändringar med ett lösenord.  
Aktivera skydd  
Markera textområde.  
Välj Infoga - Område - Skrivskydd - Skydda - Med lösenord. (Om området redan finns:  
Format - Områden.) Ange ett lösenord som består av minst 5 tecken och bekräfta det.  
Avaktivera skydd  
Välj Format - Områden - Skrivskydd, upphäv markering i rutan Skyddat.  
Ange rätt lösenord.  
Skydda celler i %PRODUCTNAME Writer-texttabell  
Innehållet i enskilda celler i en %PRODUCTNAME Writer-texttabell kan skyddas mot ändringar.  
Aktivera skydd  
Sätt markören i en cell eller markera celler.  
Välj Format - Cell - Skydda.  
Avaktivera skydd  
Sätt markören i cellen eller markera cellerna.  
Eventuellt aktiverar du först rutan Markör i skyddade områden - Tillåt under Verktyg - Alternativ - Textdokument - Formateringshjälp.  
Välj sedan Format - Cell - Upphäv skydd.  
I Navigator markerar du tabellen och väljer sedan Tabell - Upphäv skydd på snabbmenyn.  
Med tangentkombinationen Skift+Ctrl+T upphäver du skyddet för hela den aktuella tabellen eller alla markerade tabeller.  
Automatiskt skydd i kataloger  
En innehållsförteckning eller t.ex. ett sakregister som har skapats automatiskt i en %PRODUCTNAME Writer-text är automatiskt skyddat mot oavsiktliga ändringar.  
Aktivera skydd  
Sätt markören i förteckningen.  
Välj Redigera förteckning på snabbmenyn.  
Markera Skyddad mot manuella ändringar under fliken Förteckning.  
Avaktivera skydd  
Sätt markören i förteckningen.  
Eventuellt aktiverar du först rutan Markör i skyddade områden - Tillåt under Verktyg - Alternativ - Textdokument - Formateringshjälp.  
Välj Redigera förteckning på snabbmenyn.  
Markera Skyddad mot manuella ändringar under fliken Förteckning.  
I Navigator markerar du förteckningen och väljer sedan Förteckning - Upphäv skydd på snabbmenyn.  
Skydda ramar, grafik och OLE-objekt  
Många objekt kan infogas i %PRODUCTNAME -dokument.  
Du kan skydda infogad grafik efter innehåll, position och / eller storlek.  
Motsvarande gäller för ramar (i Writer) och OLE-objekt.  
Aktivera skydd  
Till exempel för ett infogat grafikobjekt i Writer: välj Format - Grafik - fliken Tillägg, området Skydda.  
Markera Innehåll, Position och / eller Storlek.  
Avaktivera skydd  
Upphäv markeringen framför någon eller några av rutorna.  
Skydda ritobjekt och formulärobjekt  
Ritobjekten som du infogar via utrullningslisten Ritfunktioner i dina dokument kan skyddas mot oavsiktlig flyttning och ändring av storleken.  
Motsvarande gäller för formulärobjekt som har infogats via utrullningslisten Formulärfunktioner.  
Aktivera skydd  
Välj Format - Position och storlek - fliken Position eller fliken Storlek.  
Markera rutan Skydda.  
Avaktivera skydd  
Välj Format - Position och storlek - fliken Position eller fliken Storlek.  
Upphäv markeringen i rutan Skydda.  
Skydda tillgång till servrar via WebDAV och FTP  
%PRODUCTNAME snabbstart i Windows  
Det finns flera möjligheter att aktivera snabbstart av %PRODUCTNAME under Windows:  
Använd kryssrutan Ladda %PRODUCTNAME vid systemstart under Verktyg - Alternativ - %PRODUCTNAME - Arbetsminne.  
Aktivera utan att starta om systemet: starta programmet quickstart.exe i katalogen {installpath }\program.  
Använd snabbstartikonen  
Om du klickar med höger musknapp på ikonen på aktivitetsfältet öppnas en undermeny.  
Här kan du bland annat öppna ett nytt tomt dokument, dialogrutan Mallar och dokument eller en Arkiv-Öppna-dialogruta.  
Om du dubbelklickar på ikonen öppnas dialogrutan Mallar och dokument.  
Kommandot Ladda %PRODUCTNAME vid systemstart kan vara aktiverat (med bock) eller inaktiverat (utan bock).  
Om det finns en bock framför kommandot och du klickar på det tas länken till quickstart.exe bort från Autostart-gruppen i Windows.  
Om det inte finns någon bock framför kommandot och du klickar på det kopieras en motsvarande länk till Autostart-gruppen.  
Kommandot Avsluta snabbstart tar bort ikonen från aktivitetsfältet och alla %PRODUCTNAME programrutiner från arbetsminnet under förutsättning att alla %PRODUCTNAME -dokument har stängts innan.  
Ta bort %PRODUCTNAME från minnet  
Stäng alla öppna %PRODUCTNAME -dokument genom att t.ex. välja Arkiv - Avsluta.  
Öppna snabbmenyn för ikonen på aktivitetsfältet.  
Välj kommandot Avsluta snabbstart.  
Nu har %PRODUCTNAME tagits bort från arbetsminnet.  
Acceptera eller ignorera ändringar  
När du får tillbaka ett dokument där andra författare har registrerat sina ändringar, kan du godta eller avslå ändringarna en och en eller alla på en gång.  
Om du har skickat ut flera kopior av dokumentet, så fogar du först samman dem till ett dokument (se ovan).  
Öppna dokumentet och välj Redigera - Ändringar - Acceptera eller ignorera....  
Dialogrutan Acceptera eller ignorera ändringar visas.  
Markera en ändring under fliken Lista i dialogrutan.  
Ändringen markeras och visas i dokumentet och du kan nu acceptera eller avböja ändringen genom att klicka på motsvarande kommandoknapp i dialogrutan.  
Om en författare har ändrat en annan författares ändring, visas detta i en hierarkisk uppställning, som du öppnar genom att klicka på plustecknet.  
Det finns även andra begränsningsalternativ.  
Du kan även filtrera efter beskrivningarna och använda platshållare (som vid reguljära uttryck i Sök och Ersätt-dialogrutan) vid inmatningen av filtret.  
I textdokument visas de ändringar som ännu inte har accepterats i listan.  
Accepterade ändringar tas bort från listan och visas i texten utan extra markering.  
På så sätt kan du även i fortsättningen se vilka ändringar som har accepterats om du vill.  
Posterna är färgkodade och informerar om resultatet av det inställda filtret.  
Svarta poster kan du acceptera eller avslå och de motsvarar filterkriterierna.  
Blåa poster motsvarar själva inte filterkriterierna, men har underordnade poster som har registrerats av filtret.  
De gröna posterna motsvarar visserligen filtret men kan ändå inte accepteras eller avslås.  
Jämföra versioner av ett dokument  
Kanske har någon av de personer som har fått en kopia av dokumentet gjort ändringar utan att registrera dem med kommandot Redigera - Ändringar - Registrera.  
Du kan antingen be personen göra om ändringarna och registrera dem i %PRODUCTNAME, eller så kan du själv jämföra kopian av dokumentet med originalet.  
Öppna originaldokumentet och välj Redigera - Jämför dokument...  
En dialogruta öppnas där du väljer kopian av dokumentet.  
Bekräfta dialogrutan.  
Nu sammanfogar %PRODUCTNAME båda versionerna i originaldokumentet.  
Alla textställen som förekommer i originaldokumentet, men inte i kopian markeras som infogade och alla ställen som saknas i originalet markeras som raderade.  
Du kan nu acceptera "infogningarna", då finns de motsvarande texterna kvar i originalet, eller acceptera "raderingarna", då infogas inte den motsvarande markerade texten, som finns i kopian, i dokumentet.  
Sammanfoga versioner  
Det är inte alltid så att ett och samma dokument ändras av olika författare och skickas vidare från en författare till nästa.  
Det är ofta bättre att ge varje författare en egen kopia av dokumentet.  
Då får du tillbaka ett antal kopior med olika ändringar i varje kopia.  
De här dokumenten kan du sedan enkelt sammanfoga i ditt originaldokument.  
Dokumenten får bara skilja sig åt när det gäller de registrerade ändringarna - för övrigt måste dokumenten vara identiska.  
Öppna originaldokumentet där du vill sammanfoga alla kopiorna igen.  
Välj Redigera - Ändringar - Sammanfoga dokument.  
En dialogruta öppnas där du väljer en kopia av dokumentet.  
Efter sammanfogningen ser du de registrerade ändringarna från kopian i originaldokumentet.  
Registrera ändringar  
Revideringsfunktionen är tillgänglig för text - och tabelldokument i %PRODUCTNAME.  
Alla typer av ändringar registreras inte (t.ex. ändring av en tabulering från vänsterjusterad till högerjusterad registreras inte).  
Men alla vanliga ändringar som en korrekturläsare gör registreras, d.v.s. kompletteringar, strykningar och ändringar av texter, vanliga formateringar och så vidare.  
1.  
Du aktiverar revideringsfunktionen genom att öppna det dokument som ska redigeras, välja Redigera - Ändringar och markera Registrera.  
2.  
Gör nu dina ändringar.  
När du skriver ny text stryks den under, medan all text som du raderar finns kvar men stryks igenom och visas i färg.  
3.  
När du placerar muspekaren på en markerad ändring visas information om typ av ändring, författaren, datum och klockslag i tipshjälpen.  
Om den aktiva hjälpen är aktiverad (på menyn Hjälp) kan du dessutom se en eventuell kommentar till ändringen.  
När du ändrar i en cell i ett tabelldokument markeras cellen med en röd kant.  
Om du sedan pekar med musen på cellen visas information om ändringen i tipshjälpen.  
Du kan förse varje markerad ändring med en kommentar genom att placera textmarkören i det ändrade området och sedan välja Redigera - Ändringar - Kommentar.  
Kommentaren visas förutom i den aktiva hjälpen också i listan i dialogrutan Acceptera eller ignorera ändringar.  
Du stänger av funktionen för registrering av ändringar genom att välja Redigera - Ändringar - Registrera på nytt.  
Bocken framför kommandot försvinner och du kan nu spara dokumentet och lämna tillbaka det till den som har bett dig om ändringarna.  
Det kan t.ex. vara ett rött streck i sidmarginalen.  
Du väljer typ av extra ändringsmarkering under Verktyg - Alternativ... - Textdokument - Ändringar eller Verktyg - Alternativ... - Tabelldokument - Ändringar.  
Här bestämmer du hur och med vilken färg som ändringarna ska markeras, var på textsidan markeringsstrecket ska vara och så vidare.  
Skydda registrering  
I ett dokument kan du registrera ändringar antingen genom att välja Redigera - Ändringar - Registrera eller Redigera - Ändringar - Skydda registrering.  
Om du har valt Skydda registrering måste du ange ett lösenord innan du kan stänga av funktionen eller acceptera eller ignorera ändringarna.  
Välj Skydda registrering.  
Dialogrutan Mata in lösenord öppnas.  
Ange ett lösenord som omfattar minst 5 tecken och bekräfta det.  
Klicka på OK.  
Versionsadministration  
På menyn Arkiv finns kommandot Versioner.  
Versionerna gör att du kan spara flera versioner av samma dokument i samma fil.  
Du kan välja att visa de enskilda versionerna eller visa skillnaderna mellan versionerna med färgmarkeringar.  
Du väljer vilka versioner av ett dokument som du vill öppna i en listruta i dialogrutan Öppna.  
Registrera och visa ändringar  
Detta gör du med revideringsfunktionen (markering av ändringar, redlining).  
När dokumentet redigeras slutgiltigt kan man gå igenom de olika ändringarna och bestämma vilka som ska tas med och vilka som ska tas bort.  
Tänk dig att du är redaktör och ska leverera ett reportage.  
Innan publiceringen läser även chefredaktören och korrekturläsaren reportaget och var och en skriver in sina ändringar.  
Chefredaktören skriver kanske "vassare formulering här" efter ett stycke och stryker ett annat helt och hållet.  
Korrekturläsaren stavningskontrollerar texten enligt gällande standard och frågar när det gäller främmande ord om du inte hellre vill använda ett svenskt uttryck.  
Du får tillbaka det redigerade dokumentet med bådas ändringsförslag och kan godta eller förkasta dem.  
Du får tillbaka kopian med kollegans kompletteringar.  
Eftersom alla kollegor och chefer arbetar med %PRODUCTNAME på ditt företag är det nu mycket enkelt att göra ett slutgiltigt dokument av resultaten.  
Skapa runda hörn  
Om du infogar en förklaring eller en rektangel med ritfunktionerna, och funktionen Redigera punkter är aktiverad, visas en liten ruta i objektets övre vänstra hörn.  
Den här ramen visar hur mycket hörnen är avrundade på objektet.  
Om den befinner sig överst till vänster blir hörnen inte avrundade; om den befinner sig på handtaget överst i mitten av objektet blir hörnen maximalt avrundade.  
Om ramen befinner sig någonstans där emellan får rundningen ett mellanliggande värde.  
Om Du för muspekaren över rutan, förvandlas den till en liten hand.  
Du kan då trycka ned musknappen och dra rutan och på så sätt ändra hörnrundningen.  
En stor kontur ger en antydan om förändringen.  
Så här skickar du ett standardfax  
Det finns två alternativ om du vill skicka ett standardfax till flera faxmottagare:  
Antingen kan du ange flera mottagare för samma dokument om faxdrivrutinen tillåter det,  
eller skicka ett dokument som ett standardbrev (kopplad utskrift) med några individuella data till var och en av mottagarna.  
Det finns mer information om standardbrev (kopplad utskrift) i %PRODUCTNAME -hjälpen.  
Tänk dock på att faxdrivrutinen måste överta den individuella tilldelningen av ett dokument till ett faxnummer.  
I allmänhet måste du skriva in en rad styrtecken och önskat faxnummer på dokumentets första rad.  
Mer information finns i dokumentationen till faxprogrammet.  
Infoga fast mellanrum, bindestreck, villkorligt skiljetecken  
Fast mellanrum  
Om du vill att ett mellanrum som ligger mellan två ord vid radslutet inte skall leda till en radbrytning, håller du ner Kommando Ctrl när du gör mellanslaget.  
Det är användbart mellan "t" och "e "(i t ex) eller mellan titeln "Dr" och personens namn.  
Skyddat bindestreck  
Ett exempel är ett företagsnamn som A-Ö.  
I det här fallet är det knappast önskvärt att A står i slutet på en rad och att Ö står i början på nästa rad.  
Tryck på Skift+Ctrl - d.v.s. håll ner skifttangenten och Ctrl-tangenten och tryck på minustangenten.  
Bindestreck, tankstreck  
Om du vill mata in längre streck använder du alternativet Ersätt tankstreck under Verktyg - AutoKorrigering / AutoFormat - Alternativ.  
Det här alternativet ersätter under vissa omständigheter ett eller två minustecken med ett längre tankstreck (se %PRODUCTNAME -hjälp).  
För andra ersättningar använder du ersättningstabellen under Verktyg - AutoKorrigering / AutoFormat - Ersättning.  
Här kan du bland annat ange att en förkortning som du bestämmer automatiskt ska ersättas av ett valfritt bindestreck vid inmatningen, t.o.m. i ett annat teckensnitt.  
Användardefinierat bindestreck  
Om du vill stödja den automatiska avstavningen genom att själv mata in bindestrecken i orden, använder du tangentkombinationen Kommando Ctrl +minustecknet.  
Ordet avstavas då på det angivna stället i radslutet även om den automatiska avstavningen inte är aktiv för det här stycket.  
Specialtecken  
Installera skrivare, fax och teckensnitt i Unix  
I Unix medföljer administrationsprogrammet för skrivare, spadmin, som hjälper dig att installera skrivare, fax och teckensnitt för %PRODUCTNAME.  
Administrationsprogrammet för skrivare, spadmin, startar du på följande sätt:  
Växla till katalogen {installpath} / program.  
Mata in:  
. / spadmin  
Efter starten ser du fönstret för administrationsprogrammet för skrivare, spadmin, där du kan göra alla viktiga inställningar.  
Vid en nätverksinstallation loggar först systemadministratör en in sig som användare root i systemet och startar administrationsprogrammet för skrivare, spadmin.  
Root-användaren skapar då en allmän skrivarkonfigurationsfil {installpath} / share / psprint / psprint.cfg för alla användare.  
Alla ändringar är direkt tillgängliga för alla användare i %PRODUCTNAME.  
Systemadministratören kan också lägga till teckensnitt för alla användare i nätverksinstallationen; men de är först tillgängliga när %PRODUCTNAME har startats om.  
Installera skrivare  
%PRODUCTNAME för Unix har bara direkt stöd för PostScript-skrivare.  
Andra skrivare måste installeras som beskrivs i avsnittet Skrivardrivrutiner i %PRODUCTNAME.  
Om du vill använda utökade egenskaper för din skrivare kan du lägga till fler skrivare.  
Lägga till skrivare  
Klicka på Ny skrivare.  
Välj alternativet Skapa en skrivare och klicka på Nästa.  
Välj en lämplig drivrutin för din skrivare.  
Om du inte använder någon PostScript-skrivare eller om din modell inte finns med, använder du drivrutinen "Generic Printer" eller så följer du beskrivningen nedan.  
Här kan du också lägga till nya drivrutiner med kommandoknappen Importera eller radera drivrutiner som inte längre behövs med kommandoknappen Radera (för mer information, se nedan).  
Sedan klickar du på Nästa.  
Markera en kommandorad med vilken det går att skriva ut på din skrivare (t.ex. lp -d my_queue).  
Klicka på Nästa.  
Ge skrivaren ett namn och bestäm om den ska vara standardskrivare.  
Klicka på Färdigställ.  
Klicka på Testsida så att en testsida skrivs ut.  
Om testsidan inte skrivs ut eller inte skrivs ut korrekt kontrollerar du alla inställningar enligt beskrivningen under Ändra skrivarinställningar.  
Från och med nu är din nya skrivare tillgänglig i %PRODUCTNAME.  
Skrivardrivrutiner i %PRODUCTNAME  
Om du installerar en icke-PostScript-skrivare måste du ställa in ditt system så att PostScript kan konverteras till skrivarens språk.  
Vi rekommenderar att du använder vanlig konverteringsprogramvara för PostScript som t.ex. Ghostscript (http: / /www.cs.wisc.edu / ~ghost /).  
I det här fallet bör du installera "Generic Printer".  
Tänk på att ställa in sidmarginalerna korrekt.  
Information om detta hittar du i de följande avsnitten.  
Om du har en PostScript-skrivare bör du alltid installera en beskrivningsfil (PostScript Printer Definition - PPD) som passar till skrivaren.  
Då kan du använda urvalet av pappersmagasin, eventuell duplexutskrift och alla installerade teckensnitt.  
Du kan också använda den generiska skrivardrivrutinen eftersom den innehåller de viktigaste uppgifterna och är lämplig för de flesta skrivare.  
I så fall måste du avstå från urvalet av pappersmagasin och ställa in sidmarginalerna rätt.  
Några PPD-filer är förinstallerade.  
Om ingen PPD-fil är installerad som är lämplig för din skrivare, hittar du olika PPD-filer under http: / /www.adobe.com / products / printerdrivers /.  
Du kan också fråga efter PPD-filer hos tillverkaren till din skrivare.  
Den lämpliga drivrutinen packar du upp med unzip och integrerar i ditt system med spadmin.  
Gör så här:  
Du kan importera eller radera drivrutiner medan du skapar en ny skrivare.  
Om du vill importera nya drivrutiner klickar du på Importera i dialogrutan med tillgängliga drivrutiner.  
Via Genomsök kan du välja ut katalogen där du har packat upp PPD-filerna.  
Klicka därefter på OK.  
Om du vill radera en skrivardrivrutin markerar du skrivardrivrutinen och klickar på kommandoknappen Radera.  
Tänk på att inte radera den generiska skrivardrivrutinen och på att raderade drivrutiner från nätverksinstallationer inte heller längre är tillgängliga för andra användare som använder samma nätverksinstallation.  
Om skrivaren har fler teckensnitt än de vanliga standardteckensnitten för PostScript, måste du även ladda AFM-filerna till dessa ytterligare teckensnitt.  
Kopiera AFM-filerna till katalogen {installpath} / share / psprint / fontmetric i %PRODUCTNAME -installationen eller till katalogen {installpath} / user / psprint / fontmetric i användarinstallationen.  
AFM-filer hittar du t.ex. på ftp: / /ftp.adobe.com / pub / adobe / type / win / all / afmfiles /.  
Ändra skrivarinställningar  
Välj skrivaren i listrutan Installerade skrivare i administrationsprogrammet för skrivare, spadmin, och klicka på Egenskaper.  
Du ser dialogrutan Egenskaper med flera flikar.  
Här kan du göra inställningarna som är tillgängliga motsvarande den valda skrivarens PPD-fil.  
Under fliken Kommando väljer du kommandot.  
Du kan ta bort överflödiga kommandon från listan genom att klicka på Ta bort.  
Under fliken Papper kan du bl.a. ange vilket pappersformat och pappersmagasin som ska användas som standard för den här skrivaren.  
Under fliken Enhet aktiverar du speciella alternativ för din skrivare.  
Om din skrivare bara kan skriva ut i svartvitt måste "Gråskalor" ställas in under Färg, annars "Färg ".  
Om omställningen till gråskalor leder till dåliga resultat kan du också välja "Färg" under Färg och överlåta omställningen åt skrivaren eller PostScript-emulatorn.  
Under den här fliken kan du också ställa in hur exakt färgerna beskrivs samt PostScript Level.  
Under fliken Teckensnittsersättning kan du välja ett skrivarteckensnitt som finns på din skrivare för varje teckensnitt som är installerat på din dator.  
På det sättet har du möjlighet att hålla nere datamängden som överförs till skrivaren.  
Teckensnittsersättningen kan aktiveras eller deaktiveras för varje skrivare.  
Om du använder den generiska skrivardrivrutinen bör du dessutom ställa in sidmarginalerna (kanten som inte kan skrivas ut) rätt under fliken Fler inställningar, så att dina utskrifter inte klipps av.  
I fältet Kommentar kan du mata in en beskrivning som också visas i dialogrutan Skriv ut.  
En del av de här inställningarna kan du också göra i dialogrutan Skriv ut eller i dialogrutan Skrivarinställningar i %PRODUCTNAME via kommandoknappen Egenskaper för varje dokument / utskrift.  
Byta namn på eller radera skrivare  
Välj en skrivare i listrutan Installerade skrivare.  
Klicka på kommandoknappen Byt namn för att byta namn på den valda skrivaren.  
Mata in ett lämpligt namn i dialogrutan som sedan visas och klicka på OK.  
Namnet måste vara entydigt och man bör kunna känna igen skrivare och användning.  
Skrivarnamn bör vara samma hos alla användare eftersom den valda skrivaren finns kvar vid utbyte av dokument om skrivaren har samma namn hos mottagaren.  
Om du vill radera den markerade skrivaren klickar du på Ta bort.  
Det går inte att ta bort standardskrivaren eller en skrivare som har skapats av systemadministratören i en nätverksinstallation med den här dialogrutan.  
Välja standardskrivare  
Om du vill göra skrivaren som är markerad i listrutan Installerade skrivare till standardskrivare dubbelklickar du på skrivarens namn eller klickar på kommandoknappen Standard.  
Integrera en faxlösning  
Om ett fungerande faxpaket som t.ex. Efax eller HylaFax är installerat på din dator, kan du också lätt skicka fax med %PRODUCTNAME.  
Klicka på Ny skrivare.  
Dialogrutan Lägg till skrivare öppnas.  
Välj Anslut en faxlösning.  
Klicka på Nästa.  
Välj om du vill använda standarddrivrutinen eller en annan skrivardrivrutin.  
Klicka på Nästa.  
Om du inte använder standarddrivrutinen, väljer du en lämplig drivrutin och klickar på Nästa.  
I följande dialogruta matar du in en kommandorad som du vill adressera faxen med.  
För varje fax som skickas ersätts "(TMP)" och "(PHONE) "i kommandoraden av en temporär fil resp. av mottagarfaxens telefonnummer.  
Om "(TMP)" förekommer i kommandoraden överförs PostScript-koden i en fil, i annat fall via standardinmatningen (d.v.s. som pipe).  
Klicka sedan på Nästa.  
Ge din nya faxskrivare ett namn och bestäm om telefonnumren som är speciellt markerade i texten (se nedan) ska tas bort från utskriften eller inte.  
Klicka på Färdigställ.  
Nu kan du skicka fax genom att skriva ut på skrivaren som just har skapats.  
I dokumentet anger du faxnumret som text.  
Du kan också mata in ett fältkommando som hämtar faxnumret från den aktuella databasen.  
Faxnumret måste i varje fall inledas med tecknen @@# och avslutas med tecknen @@.  
Ett giltig angivet nummer skulle alltså vara @@#040123456@@.  
Om de här tecknen och telefonnumret inte ska skrivas ut aktiverar du alternativet Ta bort faxnummer från utmatningen under Egenskaper under fliken Kommando.  
Om inget telefonnummer anges i dokumentet uppmanas du att ange det i en dialogruta efter utskriften.  
I %PRODUCTNAME kan du aktivera en kommandoknapp som du använder när du ska skicka till en standardfax.  
Klicka med den högra musknappen på funktionslisten, välj Synliga knappar på menyn som öppnas och aktivera Skicka standardfax på undermenyn.  
Under Verktyg - Alternativ - Textdokument - Skriv ut konfigurerar du vilken fax som används när du klickar på den här knappen.  
Tänk på att skapa ett eget utskriftsjobb för varje fax, annars får den förste mottagaren alla faxen.  
I dialogrutan Arkiv - Kopplad utskrift markerar du alltså alternativet Skrivare och sedan rutan Skapa enstaka utskriftsjobb.  
Integrera en PostScript-till-PDF-konverterare  
Om en fungerande PostScript-till-PDF-konverterare som t.ex. Ghostscript eller Adobe Acrobat Distiller( TM) är installerad på din dator, är det lätt att skapa PDF-dokument med %PRODUCTNAME.  
Klicka på Ny skrivare.  
Dialogrutan Lägg till skrivare öppnas.  
Välj Anslut en PDF-konverterare.  
Klicka på Nästa.  
Välj om du vill använda standarddrivrutinen, "Acrobat Distiller "-drivrutinen eller en annan drivrutin.  
Klicka på Nästa.  
Om du inte använder standarddrivrutinen eller "Acrobat Distiller "-drivrutinen väljer du en lämplig drivrutin och klickar på Nästa.  
I följande dialogruta matar du in en kommandorad som du vill adressera PostScript->PDF-konverteraren med.  
Dessutom anger du här katalogen där de skapade PDF-filerna ska placeras.  
Om du inte anger någon katalog används användarens hemkatalog.  
För varje skapat PDF-dokument ersätts "(TMP)" och "(OUTFILE) "i kommandoraden av en temporär fil resp. av målfilen vars namn skapas från dokumentnamnet.  
Om "(TMP)" förekommer i kommandoraden överförs PostScript-koden i en fil, i annat fall via standardinmatningen (d.v.s. som pipe).  
Om Ghostscript eller Adobe Acrobat Distiller finns i sökvägen kan du använda en av de fördefinierade kommandoraderna.  
Klicka på Nästa.  
Ge din nya PDF-konverterare ett namn.  
Klicka på Färdigställ.  
Nu kan du skapa PDF-dokument genom att skriva ut på konverteraren som just har skapats.  
Ställa in teckensnitt  
När du arbetar med %PRODUCTNAME kommer du kanske att märka att antalet teckensnitt varierar beroende på dokumenttyp.  
Det beror på att bara de teckensnitt är tillgängliga som går att använda i respektive tillämpningsfall.  
När du arbetar med ett textdokument visas bara de teckensnitt som går att skriva ut i urvalet, eftersom det är meningen att man ska kunna få ut sina dokument på papper.  
Vid ett HTML-dokument eller i onlinelayout har du bara möjlighet att använda teckensnitt som är tillgängliga på bildskärmen.  
I tabelldokument och teckningar finns däremot alla teckensnitt som antingen kan skrivas ut eller visas på bildskärmen.  
%PRODUCTNAME försöker att få visningen på bildskärmen att överensstämma med utskriften (WYSIWYG).  
Möjliga problem vid användning av teckensnitt visas vid undre kanten i dialogrutan Format - Tecken.  
Lägga till teckensnitt  
Du kan integrera ytterligare teckensnitt i %PRODUCTNAME.  
Teckensnitt som är integrerade på det här sättet är bara tillgängliga för %PRODUCTNAME och kan användas med olika Xservrar utan att de måste installeras där.  
Om du även vill göra teckensnitten tillgängliga för andra program ska du göra som vanligt; genom att lägga till teckensnitten till din Xserver. %PRODUCTNAME kan visa och skriva ut både PostScript Type1-teckensnitt och TrueType-teckensnitt (inklusive TrueType Collections).  
Om du vill integrera ytterligare teckensnitt i %PRODUCTNAME gör du så här:  
Starta spadmin.  
Klicka på kommandoknappen Teckensnitt.  
I dialogrutan som visas är alla teckensnitt som har lagts till för %PRODUCTNAME listade.  
Här kan du ta bort markerade teckensnitt med kommandoknappen Ta bort eller lägga till nya teckensnitt med kommandoknappen Lägg till.  
Klicka på kommandoknappen Lägg till.  
Dialogrutan Lägg till teckensnitt visas.  
Ange katalogen som innehåller teckensnitten som du vill lägga till.  
Klicka på... och välj ut katalogen i dialogrutan för sökvägsurval eller mata in katalogen direkt.  
Nu visas en lista över teckensnitten som finns i den här katalogen.  
Markera alla teckensnitt som du vill lägga till.  
Om du vill lägga till alla teckensnitt klickar du på kommandoknappen Markera alla.  
Med kryssrutan Skapa bara softlinks kan du bestämma om teckensnitten ska kopieras till %PRODUCTNAME -katalogen eller om bara symboliska länkar ska skapas där.  
Om teckensnitten som ska läggas till finns på ett datamedium som inte är tillgängligt hela tiden (som t.ex. en cd-rom) bör du kopiera teckensnitten.  
Klicka på kommandoknappen OK.  
Teckensnitten läggs nu till.  
Vid en nätverksinstallation installeras teckensnitten i den om möjligt.  
Om användaren inte har några skrivrättigheter här installeras teckensnitten i användarinstallationen, så att användaren som installerar dem har tillgång till dem.  
Radera teckensnitt  
Om du vill radera teckensnitt igen gör du så här:  
Starta spadmin.  
Klicka på kommandoknappen Teckensnitt.  
I dialogrutan som visas är alla teckensnitt som har lagts till för %PRODUCTNAME listade.  
Markera de teckensnitt som du vill radera och klicka på kommandoknappen Radera.  
Du kan bara radera teckensnitten som har lagts till för %PRODUCTNAME.  
Byta namn på teckensnitt  
Du kan byta namn på teckensnitt som har lagts till för %PRODUCTNAME.  
Detta är framför allt lämpligt att göra för teckensnitt som innehåller flera lokaliserade namn (som t.ex. ett engelskt och ett japanskt namn).  
Det finns även teckensnitt som innehåller ett oläsligt namn; det kan du ersätta med ett lämpligt namn.  
Starta spadmin  
Klicka på kommandoknappen Teckensnitt.  
Markera teckensnittet som du vill byta namn på och klicka sedan på kommandoknappen Byt namn.  
I dialogrutan som visas anger du ett nytt namn.  
Om teckensnittet innehåller flera namn står de som förslag i kombinationsfältet där du matar in det nya namnet.  
Klicka på OK.  
Om du markerar flera teckensnitt som du vill byta namn på visas en dialogruta för varje teckensnitt.  
Om du har valt en TrueType Collection (TTC) visas en dialogruta för varje teckensnitt som finns i den.  
Ändra standardmall  
Om du öppnar ett dokument från Arkiv-menyn - Nytt visas ett tomt dokument som baserar på en %PRODUCTNAME -standardmall, det vill säga t.ex. ett tomt text - eller tabelldokument.  
Du kan redigera och ändra det här dokumentet eller ersätta det med ett annat dokument, så att du, när du öppnar ett nytt dokument, omedelbart får upp ditt personliga dokument.  
Ändra standardmall  
Öppna först ett nytt, tomt dokument och utforma det på ett sådant sätt att det ser ut på det sätt som du vill att en mall ska se ut.  
Ändra t.ex. formatmallarna i Stylist.  
Om det redan finns ett %PRODUCTNAME -dokument som uppfyller dina krav bortfaller den här punkten naturligtvis.  
Du kan definiera dokumentmallar för alla %PRODUCTNAME -moduler.  
Nedan beskriver vi hur du definierar ett textdokument som mall.  
1.  
Spara nu dokumentet genom att välja Dokumentmall - Spara på Arkiv -menyn och t.ex. placera dokumentet i kategorin Standard.  
2.  
Välj Arkiv - Dokumentmall - Administrera  
3.  
Dubbelklicka på posten Standard i den vänstra listrutan.  
De användardefinierade dokumentmallarna i katalogen {installpath }\user\template visas.  
Markera dokumentet som du just har sparat och öppna snabbmenyn eller öppna undermenyn till kommandoknappen Kommandon.  
4.  
Välj Definiera som standardmall.  
Det är allt.  
När du öppnar ett nytt textdokument nästa gång motsvarar det nya dokumentet den mall som du har valt.  
Återställa standardmall  
Om den ändrade textmallen ska återställas till den ursprungliga standardmallen gör du så här:  
Välj Arkiv - Dokumentmall - Administrera.  
Välj snabbmenykommandot Återställ standardmall.  
På undermenyn väljer du dokumenttypen vars förinställning du vill återställa.  
När du sedan öppnar ett tomt textdokument motsvarar det återigen %PRODUCTNAME -standardmallen för textdokument.  
Så här använder du egna dokumentmallar  
Det finns några olika sätt att underlätta arbetet med egna dokumentmallar.  
En viktig punkt är göra mallarna snabbt åtkomliga.  
Du kan spara de egna mallarna på olika ställen i %PRODUCTNAME; och därför öppnar du ett nytt dokument som baserar på en av dina mallar på olika sätt.  
Mallar i mallmappen  
Du kan spara en ny mall via Arkiv - Dokumentmall - Spara eller välja filtypen "Mall" i den "normala "Spara-dialogrutan.  
När du sparar mallen i mappen {installpath} / user / template har du alltid tillgång till den via Arkiv - Nytt - Mallar och dokument.  
När du öppnar mallen skapas ett nytt namnlöst dokument som baserar på den här mallen.  
Du kan behöva uppdatera mallvyn i dialogrutan innan du kan se en ny mall.  
Välj Arkiv - Dokumentmall - Administrera och i dialogrutan väljer du Uppdatera på undermenyn till kommandoknappen Kommandon.  
Om du vill ändra mallen själv kan du öppna filen via Arkiv - Dokumentmall - Redigera och redigera den.  
Dokumentmallar  
Flytta, radera eller kopiera ikoner  
Om du vill flytta en ikon håller du ner Alternativ Alt -tangenten och drar ikonen till den nya platsen.  
När du drar en ikon till en annan plats på samma symbollist flyttas den, mellan symbollister kopieras den.  
Om du vill radera en ikon från en symbollist håller du ner Alternativ Alt -tangenten och drar ikonen till en plats där det inte finns någon list.  
Om du vill infoga eller radera det vertikala streck som finns mellan vissa ikoner eller grupper av ikoner använder du samma metod och drar en ikon lite åt sidan.  
Byta objektlister med snabbmeny  
Om markören t.ex. står i en texttabell ställs ikonerna för redigering av tabeller automatiskt till förfogande.  
Om markören står i en punktuppställning innehåller objektlisten ikoner som används till punktuppställningar.  
Om markören står i en punktuppställning i en tabell kan du byta mellan objektlisterna så här:  
Klicka på den sista ikonen på den högra sidan av objektlisten.  
Eller öppna snabbmenyn på objektlisten.  
Där finns en lista över de möjliga objektlisterna, klicka på den som du vill arbeta med.  
%PRODUCTNAME kommer ihåg vilken objektlist som du har valt i vilket sammanhang och visar den först nästa gång.  
Förbinda och dela celler  
Du kan markera celler som ligger intill varandra tillsammans och sedan sammanfoga dem till en enda cell.  
Omvänt är det möjligt att dela upp en stor cell som har sammanfogats av flera celler till enskilda celler igen.  
Kommandona är olika i %PRODUCTNAME Writer och Calc:  
Sammanfoga celler i %PRODUCTNAME Writer  
Markera de intilliggande cellerna.  
Välj Format - Cell - Förbind.  
Dela cell i %PRODUCTNAME Writer  
Placera markören i cellen som ska delas.  
Välj Format - Cell - Dela.  
I en dialogruta kan du välja om du vill dela cellen i två eller fler celler i horisontell eller vertikal riktning.  
Sammanfoga celler i %PRODUCTNAME Calc  
Markera de intilliggande cellerna.  
Välj Format - Sammanfoga celler - Definiera.  
Upphäva sammanfogade celler i %PRODUCTNAME Calc  
Placera markören i cellen som ska delas.  
Välj Format - Sammanfoga celler - Upphäv.  
Infoga och redigera tabulator  
Du sätter en tabulator genom att klicka med musen på linjalen.  
Alternativt kan du sätta tabbar i dialogrutan Format - Stycke.  
Båda sätten påverkar det aktuella stycket eller alla markerade stycken.  
Info:  
Om du vill tilldela den aktuella styckeformatmallen tabbarna, öppnar du dialogrutan Styckeformatmall (snabbmenyn till stycket, välj Redigera styckeformatmall) och matar in tabbarna där.  
Om du klickar med musen på linjalen så sätts en vänsterjusterad tabulator.  
Om du klickar med höger musknapp direkt på en tabulator på linjalen visas en snabbmeny där du kan ändra typ av tabulator.  
Om du t.ex. vill sätta flera decimaltabbar efter varandra finns det ett förenklat sätt att göra det: klicka så ofta på tabulatorsymbolen till vänster bredvid linjalen tills den önskade tabulatortypen visas och sätt tabbarna genom att klicka på linjalen.  
Urval  
Beskrivning:  
Sätta vänsterjusterad tabb  
Sätta högerjusterad tabb  
Sätta decimaltabb  
Sätta centrerad tabb  
Genom att dubbelklicka på linjalen öppnar du dialogrutan Stycke.  
Därefter visas dialogrutan Stycke med fliken Tabulator.  
Flytta tabbarna på linjalen  
En enskild tabulator flyttar du på linjalen genom att dra med musen.  
Om du vill flytta flera tabbar på linjalen trycker du på skifttangenten och håller ner den.  
Om du håller ner skifttangenten och drar en tabulator flyttas tabulatorn och alla tabbar som ligger till höger om dem.  
Avståndet mellan själva tabbarna ändras inte.  
Om du håller ner Kommando Ctrl -tangenten i stället för skifttangenten medan du drar en tabulator på linjalen, flyttas den här tabulatorn och alla tabbar som står till höger om den.  
Avstånden mellan tabbarna ändras proportionellt i förhållande till deras avstånd till sidmarginalen.  
Ändra egenskaperna för en tabulator  
När du har klickat på en tabulator på linjallisten kan du öppna dess snabbmeny och sedan ändra tabulatortypen.  
Radera en tabulator  
Du kan radera en tabulator med musen genom att dra ut den ur linjallisten samtidigt som du håller ner musknappen.  
Ändra förinställningar  
Om du vill ändra inställningen av dina standardtabbar kan du göra detta under Verktyg - Alternativ - Textdokument - Allmänt Verktyg - Alternativ - Tabelldokument - Allmänt Verktyg - Alternativ - Teckning - Allmänt Verktyg - Alternativ - Presentation - Allmänt.  
Med linjallistens snabbmeny kan du ändra den visade enheten till bl.a. centimeter, tum, punkter eller pica.  
Dessa ändringar är bara giltiga tills du avslutar %PRODUCTNAME och de gäller bara den linjal på vars snabbmeny du har gjort ändringen.  
Om du vill ändra måttenheten för linjaler permanent väljer du Verktyg - Alternativ - Textdokument - Allmänt och ändrar måttenheten där.  
Linjal  
Ändra textfärg  
Om du klickar på ikonen Teckenfärg och håller ner musknappen visas en utrullningslist där du kan välja bland fördefinierade färger.  
Teckenfärg  
Teckenfärg (andra moduler)  
Om du klickar kort på ikonen utan att någon text är markerad, ändrar muspekaren utseende och ser ut som en lutande färgburk.  
Med den här symbolen drar du över ett textområde samtidigt som du håller ner musknappen.  
Det här textområdet får då den valda färgen.  
Funktionen är aktiv så länge ikonen är "intryckt", eller tills du bara klickar utan att dra eller trycker på Esc-tangenten.  
Markera texten som ska få en annan färg och klicka sedan på den önskade färgen på utrullningslisten.  
Teckenfärg  
Växla mellan infognings - och överskrivningsläge  
Med tangentbordet:  
Tryck på Insert för att byta mellan överskrivnings - och infogningsläge.  
Det aktuella läget visas på statusraden.  
Med musen:  
Klicka på fältet med det aktuella läget (INFGA eller ÖVER) på statuslisten och växla mellan respektive läge:  
INFGA  
Infogningsläget är aktiverat.  
Textmarkören är ett blinkande lodrätt streck.  
Klicka med musen i fältet för att aktivera överskrivningsläget.  
ÖVER  
Överskrivningsläget är aktiverat.  
Textmarkören är ett blinkande block.  
Klicka med musen i fältet för att aktivera infogningsläget.  
Tangentkommandon  
Komplettering av filnamn (AutoComplete)  
Namn på kataloger och mappar kompletteras resp. skrivs in automatiskt i URL-fältet och i dialogrutorna för att öppna och spara filer så snart du trycker på tangenten Pil upp eller Pil ned.  
Om du precis har öppnat dokumentet "Brev1.sdw" från din dokumentmapp C:\Docs ser du följande URL i URL-fältet: "file: / //C_BAR_ / Docs / Brev1.sxw ".  
Om du nu dessutom vill öppna dokumentet "Brev till företaget XYZ beträffande de nya avtalen.sxw" som finns i samma mapp gör du på följande sätt:  
Klicka på URL-fältet.  
Det markeras i sin helhet.  
Tryck på den högra piltangenten.  
På det sättet avmarkeras hela URL-fältet och markören placeras i slutet av posten.  
Radera så många tecken med backstegstangenten att bara början av det nya filnamnet är kvar.  
I det här exemplet raderar du de sista tecknen i filnamnet "Brev1.sdw", så att bara "Brev" blir kvar.  
Tryck nu på Pil nedåt. %PRODUCTNAME visar nästa fil vars namn börjar med "Brev".  
Så snart den önskade filen visas trycker du på returtangenten.  
Så snart du trycker på returtangenten byts det aktuella dokumentet ut mot det nya.  
Om du vill öppna det nya dokumentet utan att stänga det gamla, trycker du på Kommando Ctrl och Retur.  
När kombinationsfältet Ladda URL i funktionslisten har markerats i sin helhet kan du bläddra genom listan på de redan markerade URL:erna med piltangenterna Pil upp och Pil ned.  
Genom att trycka på returtangenten eller Kommando Ctrl och Retur öppnar du det dokument som visas i kombinationsfältet från hårddisken eller från Internet.  
Med tangenterna PageUp och PageDown visar du det första respektive sista dokumentet i listan.  
När du har öppnat en fil med kombinationsfältet Ladda URL måste du alltså tänka på att du först måste placera markören i dokumentet med musen, innan du börjar bläddra i det med PageUp och PageDown.  
I stället för musen kan du också använda tangenten Esc för att åter placera markören i dokumentet.  
Om hela URL:en är markerad trycker du två gånger på Esc, i annat fall bara en gång.  
Om du inte klickar med musen eller trycker på Esc, bläddrar du nämligen genom posterna i kombinationsfältet.  
Öppna filer snabbt utan dialogruta  
Om du har öppnat en fil och vill öppna en till från samma mapp, och filens namn bara marginellt skiljer sig från den aktuella filens namn, kan du snabbt öppna den nya filen med hjälp av kombinationsfältet Ladda URL på funktionslisten.  
Klicka på kombinationsfältet Ladda URL till vänster i funktionslisten.  
Det innebär att du omedelbart kan skriva ett nytt namn som ersätter det gamla namnet i fältet.  
Eller så flyttar du markören med piltangenterna och redigerar det befintliga namnet.  
Om du trycker på returtangenten ersätts det aktuella dokumentet med dokumentet som nämns i URL:n.  
Om du håller ner Ctrl-tangenten när du trycker på Retur öppnas dokumentet som nämns i URL:n men det ersätter inte det aktuella dokumentet.  
Version och buildnummer, medarbetarlista  
Välj Hjälp - Om %PRODUCTNAME.  
Du ser en dialogruta med information.  
Du får mer information om du håller ner Kommando Ctrl -tangenten i den här dialogrutan och trycker på tangenterna S D T efter varandra.  
Alldeles i början visas information om versionen och buildnummer.  
Du avslutar informationen genom att trycka på returtangenten Esc-tangenten.  
OpenOffice.org  
Ändra arbetskatalog  
Om du öppnar dialogrutan för att öppna ett dokument i %PRODUCTNAME, ser du först din arbetskatalog där.  
Du kan ändra vilken katalog %PRODUCTNAME visar här på följande sätt:  
Välj Verktyg - Alternativ - %PRODUCTNAME - Sökvägar.  
Dubbelklicka på posten Arbetskatalog.  
I dialogrutan Välj ut sökväg väljer du katalogen som du vill använda som arbetskatalog och klickar på Välj ut.  
Avsluta den andra dialogrutan med OK.  
Du gör ungefär likadant när du byter ut katalogen som %PRODUCTNAME visar när du ska infoga ett grafikobjekt: ändra sökvägen för posten Grafik.  
Sökvägar  
Hjälp  
Via hjälpmenyn kan du öppna och kontrollera hjälpsystemet i %PRODUCTNAME.  
Innehåll  
Här öppnar du huvudsidan i %PRODUCTNAME -hjälpen för det aktiva programmet.  
Du kan bläddra i hjälpen efter ämne och söka efter indexord eller fri text.  
Help Agent  
Under Verktyg - Alternativ - %PRODUCTNAME - Allmänt finns en kryssruta som har samma effekt.  
Tips  
Här aktiverar och inaktiverar du visningen av tipshjälpen.  
Om tipshjälpen är aktiv visas namnet på ett element på bildskärmen när muspekaren är placerad där.  
Aktiv hjälp  
Här sätter du på och stänger av visningen av den aktiva hjälpen.  
Om den aktiva hjälpen är på visas en kort funktionsbeskrivning för ett element på bildskärmen när muspekaren är placerad där.  
Om %PRODUCTNAME  
Med det här kommandot visar du allmän information om programmet.  
Det gäller t.ex. versionsnumret och copyright.  
Funktionslist  
Funktionslisten är den översta symbollisten i %PRODUCTNAME -fönstret.  
Här finns ikoner för de viktigaste funktionerna som alltid är tillgängliga.  
Om några ikoner inte gäller i det aktuella sammanhanget gråmarkeras de och kan inte aktiveras.  
Om t.ex. ett grafikobjekt är markerat, kan ikonen Infoga tabell inte aktiveras eftersom det inte går att infoga en tabell i ett grafikobjekt.  
Dokumenttypen som skapas med enkelt musklick beror på den senast skapade dokumenttypen och representeras av den visade ikonen.  
Öppna fil  
Statuslist vid %PRODUCTNAME Basic-dokument  
Statuslisten visar information om det för tillfället öppnade %PRODUCTNAME Basic-dokumentet.  
Statuslisten kan konfigureras (under Verktyg - Anpassa).  
I normala fall ser du fält som har följande betydelse från vänster till höger:  
Hyperlänklist  
På hyperlänklisten kan du ange sökord och söka på Internet med de förinställda sökmotorerna genom att klicka med musen.  
Här kan du dessutom redigera hyperlänkar till andra dokument eller Internet.  
Du öppnar hyperlänklisten via Visa - Symbollister - Hyperlänklist.  
Databaslist  
I datakällvyn visas databaslisten i den övre kanten.  
Originaltabellen ändras inte.  
Resultatet av en sortering eller filtrering sparas automatiskt och finns kvar tills du ändrar eller ångrar sorteringen eller filtreringen.  
Om ett filter är aktivt är ikonen Använd filter på databaslisten intryckt.  
Data i text Data i text  
Kopplad utskrift  
Den här ikonen öppnar dialogrutan Kopplad utskrift.  
Här hittar du alla funktioner för att skriva ut och spara kopplade utskrifter.  
Formulärlist  
Formulärlisten i formulärvyn innehåller olika funktioner för redigering av databastabeller och styrning av datavisningen.  
Den hjälper dig att navigera i dataposterna och att infoga eller radera dataposter.  
Om en datapost sparas i formuläret, överförs ändringarna till databasen.  
Vidare innehåller formulärlisten funktioner för sortering och filtrering av data och möjliggör även olika metoder för sökning i dataposterna.  
Formulärlisten är bara synlig för formulär med databaskoppling.  
I formulärets utkastläge är den dold.  
Se även databaslisten.  
Originaltabellen ändras inte.  
En sortering eller filtrering sparas i dokumentet tills du upphäver den.  
Om ett filter har använts för formuläret är ikonen Använd filter på formulärlisten i intryckt läge.  
Du kan också ställa in sorteringar eller filtreringar i dokumentet via formuläregenskaperna (se Formuläregenskaper - fliken Data - Egenskaper Sortering och Filter).  
Om formuläret baseras på en SQL-sats (se Formuläregenskaper - fliken Data - egenskap Datakälla), är filtrerings - och sorteringsfunktionerna bara tillgängliga om den här SQL-satsen enbart refererar till en tabell och det dessutom inte är skrivet i databasens Native-SQL.  
Datapostnummer  
Här visas vilken datapost som är markerad för tillfället.  
Du kan ange ett nummer för att gå direkt till motsvarande datapost.  
Första datapost  
Med den här ikonen går Du till den första dataposten.  
Föregående datapost  
Med den här ikonen går Du till föregående datapost.  
Nästa datapost  
Med den här ikonen går Du till nästa datapost.  
Sista datapost  
Med den här ikonen går Du till den sista dataposten.  
Spara datapost  
Här sparas en ny inmatning av data och ändringarna förs in i databasen.  
Ångra: inmatning av data  
Här kan du ångra en inmatning.  
Ny datapost  
Klicka på den här ikonen om Du vill mata in en ny datapost.  
Radera datapost  
Om Du klickar på den här ikonen raderas den för tillfället markerade dataposten.  
Du måste bekräfta raderingen innan den utförs.  
Sök datapost...  
Sortera...  
SQL-sökningslist  
Om du skapar eller redigerar en sökning i sökningsutkastet kan du använda ikonerna på SQL-sökningslisten för att generera sökningen.  
Beroende på om sökningen skapas under Utkast-fliken eller SQL-fliken visas följande ikoner:  
Lägg till tabeller  
Under fliken SQL visas följande ikon:  
Objektlist för formulärutkast  
Den här objektlisten visas när ett formulär är öppet i utkastläge och du har markerat ett formulärobjekt.  
Lägg till fält  
Gruppering  
Upphäv gruppering  
Gå in i gruppering  
Lämna gruppering  
Visa raster  
Fäst mot raster  
Om du aktiverar den här ikonen, kan objekten bara flyttas mellan de olika rasterpunkterna.  
Hjälplinjer vid förflyttning  
Bézierobjektlist  
Bézierobjektlisten visas när du har markerat ett bézierobjekt och klickat på kommandot Redigera punkter.  
Här finns olika funktioner för att redigera punkter i en kurva eller ett objekt som har omvandlats till en kurva.  
Följande ikoner är tillgängliga:  
Redigera punkter  
Med ikonen Redigera punkter kan du sätta på eller stänga av redigeringsläget för bézierobjekt.  
I redigeringsläget kan enskilda punkter i ett ritobjekt markeras.  
Redigera punkter  
Flytta punkter  
När den här ikonen är aktiverad kan du flytta punkter.  
När du pekar på en av punkterna visar markören en liten tom kvadrat.  
Tryck nu ned musknappen och dra punkten till ett annat ställe.  
Kurvan på båda sidor om punkten följer rörelsen och kurvan formas om fram till nästa punkt i båda riktningar.  
Om du pekar på kurvan mellan två punkter eller på ytan i en sluten kurva, trycker ned musknappen och drar, så flyttas hela kurvan utan att formen ändras.  
Flytta punkter  
Infoga punkter  
Genom att klicka på ikonen aktiverar du infogningsläget, där du kan infoga nya punkter.  
I det här läget kan du även flytta punkter, precis som i flyttningsläget.  
Men om du klickar på kurvan mellan två punkter och flyttar musen en bit där med nertryckt musknapp, infogar du en ny punkt där.  
Punkten är en jämn punkt, linjerna till kontrollpunkterna är alltså parallella och förblir parallella även när de flyttas.  
Om Du vill skapa en hörnpunkt måste Du först infoga en jämn punkt eller symmetrisk punkt och sedan omvandla den till en hörnpunkt med ikonen Sätt hörnpunkt.  
Du kan även infoga punkter utanför den befintliga kurvan.  
Klicka i närheten av kurvan i infogningsläge så bedömer programmet automatiskt med hjälp av avstånden, mellan vilka två punkter på kurvan den nya punkten ska infogas.  
Om placeringen bedöms vara rimlig infogas den nya punkten och kurvan anpassas.  
Om Du håller Kommandotangenten Ctrl-tangenten nedtryckt när Du klickar utanför kurvan så skapar Du ett nytt kurvsegement, som inte är direkt förbundet med den befintliga kurvan.  
Men det är en kombination med den aktuella kurvan och flyttas, kopieras, raderas etc. tillsammans med den.  
Infoga punkter  
Radera punkter  
Med den här ikonen kan du radera en eller flera markerade punkter.  
Om du vill markera flera punkter håller du ner skifttangenten när du klickar på dem.  
Markera punkterna först och klicka sedan på den här ikonen.  
Du kan även trycka på Delete-tangenten.  
Radera punkter  
Dela kurvan  
Med den här ikonen delar du en kurva.  
Markera den eller de punkter där kurvan ska delas och klicka sedan på den här ikonen.  
Dela kurvan  
Omvandla till kurva  
Med den här ikonen omvandlar du en rundad kurva till en rät linje och omvänt.  
Om två punkter är markerade omvandlas kurvsegmentet mellan dem.  
Om du har markerat mer än två punkter omvandlas en annan del av kurvan varje gång du klickar på den här ikonen.  
Vid behov kan även rundade punkter omvandlas till hörnpunkter och omvänt.  
De kan inte omvandlas till rundade punkter om Du inte först omvandlar den räta linjen till en kurva igen.  
Omvandla till kurva  
Sätt hörnpunkt  
Med den här ikonen omvandlar du den aktuella punkten eller de markerade punkterna till hörnpunkter.  
Kurvan löper inte jämnt genom en hörnpunkt utan har ett hörn.  
Sätt hörnpunkt  
Jämn övergång  
Klicka på den här ikonen för att göra om en hörnpunkt eller en symmetrisk punkt till en jämn punkt.  
De båda linjerna till hörnpunktens kontrollpunkter justeras parallellt och kan bara flyttas tillsammans.  
Men linjerna till kontrollpunkterna får vara olika långa, vilket leder till olika kraftig böjning av kurvan.  
Jämn övergång  
Symmetrisk övergång  
Med den här ikonen blir en hörnpunkt eller jämn punkt till en symmetrisk punkt.  
Linjerna till kontrollpunkterna är parallellt justerade och lika långa.  
Kurvans böjning är lika kraftig åt båda hållen i en symmetrisk punkt.  
Symmetrisk övergång  
Slut Bézier  
Med den här ikonen kan du sluta den aktuella linjen.  
En linje sluts alltid genom att den sista punkten (som visas som en något förstorad kvadrat) förbinds med startpunkten.  
Detta sista delsegment av linjen öppnas alltid direkt framför startpunkten, där en ny ändpunkt infogas.  
Slut Bézier  
Reducera punkter  
Med den här ikonen märker du den aktuella punkten eller de markerade punkterna för radering.  
Detta görs om punkten ligger på en rät linje.  
Om du omvandlar en kurva eller polygon till en rät linje med ikonen Omvandla till kurva eller ändrar en kurva med musen så att den här punkten ligger på en rät linje, tas punkten bort.  
Den vinkel där punktreduktionen ska börja, ställer du in under Verktyg - Alternativ - Teckning - Raster. ställer du in under Verktyg - Alternativ - Presentation - Raster. är förinställd till 15°.  
Reducera punkter  
Mer information om datakällor i %PRODUCTNAME  
I det här avsnittet hittar du mer information om hur du arbetar med datakällor i %PRODUCTNAME.  
Registrering av systemadressboken  
Åtkomst till data i text - eller tabelldokument  
Databasfunktioner i %PRODUCTNAME  
Här finns en allmän introduktion av databaskonceptet i %PRODUCTNAME och anvisningar om hur nya datakällor ställs in och hur datakällor redigeras, hur externa datakällor används som adressbok när standardbrev (kopplad utskrift) skapas, hur databastabeller och sökningar skapas och redigeras, hur formulär skapas och hur dokument länkas till datakällor.  
Kortkommandon  
Det här avsnittet innehåller de kortkommandon som är viktiga när du använder %PRODUCTNAME.  
Facktermer enkelt förklarade (ordlista)  
I det här avsnittet hittar du en allmän ordlista över facktermerna i %PRODUCTNAME och en särskild förteckning över Internettermer.  
Programmering av %PRODUCTNAME %PRODUCTVERSION  
%PRODUCTNAME %PRODUCTVERSION kan styras med hjälp av %PRODUCTNAME API.  
%PRODUCTNAME %PRODUCTVERSION har ett nytt gränssnitt, Application Program Interface (API), som gör det möjligt att styra %PRODUCTNAME -komponenter via olika programmeringsspråk.  
Det finns ett %PRODUCTNAME %PRODUCTVERSION Development Kit till det nya programmeringsgränssnittet.  
Mer information om %PRODUCTNAME API-referens (http: / /api.openoffice.org /)  
Makron som du har skapat med %PRODUCTNAME Basic och som baserar på det gamla programmeringsgränssnittet, stöds inte längre av den aktuella versionen.  
Om du vill veta mer om %PRODUCTNAME Basic väljer du "Hjälp till %PRODUCTNAME Basic" i kombinationsfältet.  
Java  
%PRODUCTNAME stöder Java.  
Du kan köra tillämpningar, appletprogram och JavaBeans i %PRODUCTNAME.  
Nedan följer de olika avsnitten om Java som finns i %PRODUCTNAME -hjälpen.  
Om Java ska kunna fungera i %PRODUCTNAME, måste Java 2 Runtime Environment från Sun Microsystems vara installerat.  
När du installerade %PRODUCTNAME erbjöds du automatiskt att installera dessa filer, om de inte redan var installerade.  
Det är möjligt att installera filerna i efterhand.  
Den körbara setup-filen finns i %PRODUCTNAME / program-mappen och på %PRODUCTNAME -cd:n.  
I andra operativsystem eller för andra versioner ändras namnet på motsvarande sätt.  
Du måste ha aktiverat Java i %PRODUCTNAME, för att kunna köra Java-tillämpningar.  
Java aktiverar du under Verktyg - Alternativ - %PRODUCTNAME - Säkerhet.  
Ändringarna under Verktyg - Alternativ - %PRODUCTNAME - Säkerhet övertas, även om Java Virtual Machine (JVM) redan har startats.  
Även ändringarna under Verktyg - Alternativ - Internet - Proxy övertas när JVM har startats.  
Här utvärderas bara de båda raderna "Http Proxy" och "Ftp Proxy "med sina portar.  
%PRODUCTNAME och Internet  
Här hittar du information om "Internet".  
I den allmänna Internet-ordlistan förklaras de viktigaste termerna.  
Alternativ  
Det här kommandot öppnar en dialogruta för individuell anpassning av programmet.  
Ändringarna sparas automatiskt.  
Du visar innehållet under en överskrift i denna hierarkiska vy genom att klicka på plustecknet eller dubbelklicka på överskriften, och döljer det igen genom att klicka på minustecknet framför överskriften.  
När du öppnar menyn Verktyg - Alternativ för första gången visas Användardata.  
Varje gång därefter visas den senast aktiva sidan.  
Välj det område vars förinställningar du vill se eller ändra.  
%PRODUCTNAME  
Ladda / spara  
Språkinställningar  
Internet  
Textdokument  
HTML-dokument  
Tabelldokument  
Presentation  
Teckning  
Formel  
Diagram  
Datakällor  
Alternativ %PRODUCTNAME  
Här gör du allmänna inställningar för ditt arbete med %PRODUCTNAME.  
I dialogrutan ställer du bland annat in dina användardata, minne, utskrift, sökvägar till viktiga filer och kataloger och färger.  
De här inställningarna sparas automatiskt så att de alltid gäller.  
Användardata  
Här har du möjlighet att ange eller ändra olika användardata.  
De uppgifter som visas här och som du kan redigera, har du eventuellt redan angett vid installationen av %PRODUCTNAME.  
Nästan alla data används i olika mallar och av AutoPiloter i %PRODUCTNAME så att de automatiskt skrivs in i respektive fältkommandon.  
Uppgifterna i datafälten "Förnamn" och "Efternamn "används under Arkiv - Egenskaper för att t.ex. ange ditt namn som författare till ett nytt dokument.  
Användaruppgifterna Företag, Efternamn, Gata, Postadress, Titel och Befattning förs automatiskt in i en intern ordlista, så att de känns igen som rättskrivna vid rättstavningskontroll.  
Vid framtida skrivfel kan uppgifterna användas som korrigeringsförslag.  
Ändringar av uppgifterna träder i kraft först när du har startat om %PRODUCTNAME.  
Adress  
I området Adress anger eller ändrar du dina personliga användardata.  
Företag  
I det här datafältet anger du namnet på ditt företag.  
Förnamn  
Ange förnamnet här.  
Efternamn  
Ange efternamnet här.  
Initialer  
Här anger du dina initialer.  
Gatuadress  
I det här datafältet kan du ange eller ändra din gatuadress.  
Postnr / Ort  
Här anger eller ändrar du ditt postnummer.  
Ort  
Ange orten här.  
Land  
Ange i vilket land du bor.  
Titel  
Ange din titel här.  
Befattning  
Här anger du din befattning på företaget.  
Tfn (priv.)  
Ange ditt privata telefonnummer.  
Tfn. (arb.)  
Här anger du ditt telefonnummer på arbetsplatsen.  
Fax  
Här anger du ditt faxnummer.  
E-post  
Här anger du din e-postadress.  
Skriv adressen enligt mönstret "mitt.namn@min.leverantör.se" (utan citattecknen).  
Spara  
Här kan du bland annat definiera olika förinställningar som gäller när du sparar dokument samt välja standardfilformat.  
Ladda  
Ladda användarspecifika inställningar med dokumentet  
Markera den här rutan om de användarspecifika inställningar som har sparats i ett dokument ska laddas med dokumentet.  
Om rutan inte är markerad laddas inte följande information som dokumentet alltid innehåller, d.v.s. dina egna inställningar fortsätter att gälla för det här dokumentet:  
Inställningar som finns under Arkiv - Skriv ut - Fler,  
namn på faxskrivaren,  
avståndsalternativ för stycken före texttabeller,  
information om automatisk uppdatering för länkar, fältfunktioner och diagram,  
information om asiatiska teckenformateringar.  
Det finns några inställningar som alltid laddas med ett dokument, oberoende av den här kryssrutan:  
Skrivarnamn,  
datakälla som är kopplad till dokumentet och datakällans vy.  
Spara  
Redigera egenskaper innan  
Om du markerar den här rutan visas först dialogrutan Egenskaper varje gång du använder funktionen Spara som.  
Skapa alltid säkerhetskopia  
Varje gång du sparar sparas dessutom en kopia av filen med samma namn och tillägget BAK i Backup-katalogen.  
Säkerhetskopian arkiveras i den mapp som du har valt som mapp för säkerhetskopior under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar.  
I förinställningen är det mappen "Backup" i %PRODUCTNAME -user-mappen.  
Spara automatiskt var  
Om den här rutan är markerad sparar %PRODUCTNAME det aktuella dokumentet med ett tidsintervall som du har definierat, som om du hade tryckt på Ctrl+S.  
minut  
Här kan du bestämma tidsintervallet i minuter för hur ofta dokumentet ska sparas automatiskt.  
Bekräfta före spara  
Om du markerar rutan Bekräfta före spara visas en säkerhetskontroll innan dokumentet sparas automatiskt.  
Storleksoptimering för XML-format (utan pretty printing)  
Om den här rutan är markerad skriver %PRODUCTNAME XML-data utan indrag och radbrytningar när ett dokument sparas.  
Då går det snabbare att spara och öppna dokumentet och filstorleken minskar.  
Avmarkera rutan om du vill läsa XML-filer i en textredigerare med strukturerat skrivsätt.  
Spara URL:er relativt  
Här väljer du förinställningen till relativ adressering av URL:er i filsystemet och på Internet.  
Relativ adressering är bara möjlig om utgångsdokument och dokumentet, som det hänvisas till med en hyperlänk, finns på samma enhet.  
En relativ adress utgår alltid från den aktuella katalogen där det aktuella dokumentet står.  
Den absoluta adresseringen utgår däremot alltid från rotkatalogen.  
Ditt dokument finns t.ex. i katalogen / work / docs C:\work\docs.  
Dessutom finns det en katalog / work / images C:\work\images.  
Du refererar till en bild i katalogen / work / images C:\work\images på följande sätt:  
Exempel  
Filsystem  
Internet  
relativt  
.. / images / img.jpg  
.. / images / img.jpg  
absolut  
file: / //c _BAR_ / work / images / img.jpg  
http: / /myserver.com / work / images / img.jpg  
Visningen i tipshjälpen visar alltid en absolut sökväg.  
Men när du sparar i HTML-filformat anges en relativ sökväg i %PRODUCTNAME om du aktiverar det här alternativet.  
i filsystem  
Här kan du välja att URL:er ska sparas relativt i filsystemet.  
på Internet  
Här kan du väljer att URL:er ska sparas relativt på Internet.  
Standardfilformat  
Välj här vilket filformat som ska vara standard när du sparar olika dokumenttyper.  
Dokumenttyp  
Välj dokumenttypen som du vill definiera standardfilformatet för.  
Spara alltid som  
Välj filformat här.  
Dokument av typen som har valts till vänster sparas alltid i det här filformatet, såvida du inte väljer ett annat filformat i dialogrutan Spara som.  
Sökvägar  
Här definierar du sökvägarna till viktiga mappar.  
Under posten Arbetskatalog väljer du den mapp som ska visas först i dialogrutan Öppna när du öppnar ett dokument.  
På motsvarande sätt väljer du den mapp som ska visas när ett grafikobjekt öppnas under Grafik.  
Posterna för Standardmallar och AutoPilot namnger de mappar där länkarna, filerna och mapparna finns som visas som undermeny under menyerna Arkiv - Nytt och Arkiv - AutoPilot.  
Där kan du välja sökvägar till olika mappar där dina AutoTexter finns, t.ex. privata och arbetsrelaterade.  
Motsvarande gäller för posten Dokumentmallar.  
Men den kan även innehållera flera sökvägar.  
Via kommandoknapparna Redigera... - Lägg till... kan du också ange ytterligare sökvägar som ska läggas till.  
De visas åtskilda med ett semikolon.  
Du kan använda några variabler: $(inst) står för sökvägen till mappen där %PRODUCTNAME har installerats. $(user) står för den sökväg där användaren har installerat sina %PRODUCTNAME -filer under den användardefinierade installationen.  
Även sökvägsvariabeln för operativsystemet kan utläsas.  
Den heter $(path).  
Typ / Sökväg  
Om du vill ändra en av posterna i den här listrutan, markerar du den först och klickar sedan på Redigera.  
Alternativt kan du dubbelklicka på posten.  
Standard  
Den här kommandoknappen återställer de förinställda sökvägarna för alla markerade poster.  
Redigera...  
Genom att klicka en gång på den här kommandoknappen visas beroende på typ någon av dialogrutorna Välj ut sökväg eller Välj sökvägar.  
Posterna i listrutan Sökväg  
Du kan ändra posternas ordningsföljd genom att klicka på Typ.  
Kolumnbredden ändrar du genom att flytta linjen mellan kolumnerna med musen.  
I beteckningen av sökvägar står {netinstall} för %PRODUCTNAME -katalogen på nätverksservern, från vilken den enskilde användaren har utfört sin användardefinierade installation.  
Användaren har installerat i sin hemkatalog på sin hårddisk och katalogen som har skapats för %PRODUCTNAME -filerna där kallas för {userinstall}.  
Poster i listrutan Sökväg som har mer än en sökvägsangivelse  
Posterna AutoKorrigering, AutoText, Basic, Dokumentmallar samt Gallery kan innehålla mer än en sökvägsangivelse.  
I en nätverksmiljö står t.ex. några filer i katalogen {netinstall}.  
Där är de tillgängliga för alla användare men kan i vanliga fall inte ändras eftersom användarna bara har läsrättigheter där.  
AutoText-block som användaren definierar själv skapas t.ex. automatiskt i katalogen under {userinstall} där användaren även har skrivrättigheter.  
Namn  
Förinställning  
Betydelse  
Add-ins  
{netinstall} / program / addin C:\{installpath }\program\addin  
I den här mappen arkiveras alla add-ins.  
Arbetskatalog  
Standardokumentmapp i ditt system  
Den här mappen visas när du öppnar dialogrutan Öppna eller Spara.  
AutoKorrigering  
{userinstall} / user / autocorr ;{netinstall} / share / autocorr C:\{installpath}\user\autocorr; C:\{installpath }\share\autocorr  
Här sparas förinställningarna till dialogrutan AutoKorrigering.  
AutoText  
{userinstall} / user / autotext ;{netinstall} / share / autotext / swedish C:\{installpath}\user\autotext; C:\{installpath }\share\autotext / swedish  
I mapparna som nämns här arkiveras dina AutoText-block.  
BASIC  
{userinstall} / user / basic ;{netinstall} / share / basic C:\{installpath}\share\basic; C:\{installpath }\user\basic  
Här finns de %PRODUCTNAME Basic-filer som bl.a. behövs till AutoPiloterna.  
Användarkonfiguration  
{userinstall} / user / config C:\{installpath }\user\config  
Mapp för användarinställningar  
Användarordlistor  
{userinstall} / user / wordbook C:\{installpath }\user\wordbook  
Här finns de användarordlistor som du har skapat.  
Dokumentmallar  
{netinstall} / share / template / swedish ;{userinstall} / user / template C:\{installpath}\share\template\swedish; C:\{installpath }\user\template  
Mallarna kommer från de mappar och underordnade mappar som finns här.  
Filter  
{netinstall} / program / filter C:\{installpath }\program\filter  
I den här mappen finns alla filter.  
Gallery  
{netinstall} / share / gallery ;{userinstall} / user / gallery C:\{installpath}\share\gallery; C:\{installpath }\user\gallery  
Den här mappen innehåller Gallery.  
Grafik  
{netinstall} / share / gallery C:\{installpath }\share\gallery  
Den här mappen visas när du öppnar dialogrutan för att öppna eller spara ett grafikobjekt.  
Hjälpfiler  
{netinstall} / help C:\{installpath }\help  
Sökvägen till hjälpen  
Konfiguration  
{netinstall} / share / config C:\{installpath}\share\config C:\{installpath }\share\config  
Här finns konfigurationsfilerna.  
Den här posten kan inte ändras.  
Lingvistik  
{netinstall} / share / dict C:\{installpath }\share\dict  
Här arkiveras de filer som rättstavningskontrollen behöver.  
Moduler  
{netinstall} / program C:\{installpath }\program  
Här står sökvägen till modulerna.  
Standardposten ska inte ändras men Du kan lägga till ytterligare sökvägar.  
Meddelandelager  
{userinstall} / user / store C:\{installpath }\user\store  
Här lagras utgående e-post.  
Paletter  
{userinstall} / user / config C:\{installpath }\user\config  
Här står sökvägen till palettfilerna som bl.a. innehåller dina definitioner av färger, mönster och så vidare.  
Plug-ins-katalog  
{userinstall} / user / plugin ;{netinstall} / share / plugin C:\{installpath}\share\plugin; C:\{installpath }\user\plugin  
Här arkiveras plug-ins.  
Säkerhetskopior  
{userinstall} / user / backup C:\{installpath }\user\backup  
Här arkiveras de säkerhetskopior av dokument som har skapats automatiskt.  
Ikoner  
{netinstall} / share / config / symbol C:\{installpath }\share\config\symbol  
Från den här katalogen hämtas ikonerna på symbollisterna.  
Temporär baskatalog  
{userinstall} / user / temp C:\{installpath }\user\temp  
Här skapar %PRODUCTNAME sina temporära filer.  
Ordlistor  
{netinstall} / share / wordbook / swedish C:\{installpath }\share\wordbook  
Här arkiveras ordböckerna som ingår.  
Katalogstrukturen för %PRODUCTNAME  
I %PRODUCTNAME har bl.a. följande mappar och filer en särskild betydelse.  
Katalog / fil  
Betydelse  
(Din Windowsmapp för egna inställningar) - sversion.ini .sversionrc i hemkatalogen  
Den här filen identifierar den %PRODUCTNAME -version som för närvarande används.  
{installpath} / user / autotext  
Här hittar du AutoTexter som filer.  
Om du vill behålla dina autotexter måste du spara de här filerna innan du gör en ny installation.  
Se AutoText.  
{installpath} / user / backup  
Till den här katalogen säkerhetskopieras Dina dokument automatiskt, om Du har aktiverat den här funktionen.  
Se Säkerhetskopia.  
{installpath} / user / wordbook  
I den här mappen finns de ordböcker som Du har skapat för rättstavningskontrollen.  
{installpath} / share / plugin eller user / plugin  
Därför behöver du normalt sett inte installera plug-ins i den här mappen.  
Välj sökvägar / filer  
Här väljer du de mappar som innehåller AutoText-moduler eller dokumentmallar som du bör ha tillgång till i %PRODUCTNAME.  
När du ska skicka standardbrev per e-post (mailing) väljer du filerna som du vill bifoga e-breven här.  
Sökvägar / Filer  
Här visas sökvägarna eller filerna som redan har lagts till.  
Lägg till...  
Öppnar dialogrutan Välj ut sökväg där du kan välja ytterligare en mapp eller dialogrutan Öppna där du kan välja ytterligare en fil.  
Lingvistik  
Här väljer du egenskaperna för rättstavningskontroll, avstavning och synonymordlista.  
En del av de här funktionerna finns även i dialogrutan Lingvistik som du kan öppna under rättstavningskontrollen.  
Tillgängliga språkmoduler  
Här ser du vilka språkmoduler som är installerade.  
En språkmodul kan innehålla en, två eller tre underordnade moduler: rättskrivning, avstavning och synonymordlista.  
Varje underordnad modul kan finnas på en eller flera språk.  
Om du klickar framför namnet på modulen för att sätta en markering aktiverar du samtidigt alla underordnade moduler.  
Om du tar bort en markering deaktiverar du samtidigt alla underordnade moduler.  
Om du bara vill aktivera eller deaktivera enstaka underordnade moduler växlar du till dialogrutan Redigera moduler.  
Redigera  
Om du vill redigera en språkmodul markerar du en språkmodul och klicka på Redigera.  
Dialogrutan Redigera moduler visas.  
Användarordlistor  
I den här listrutan listas de tillgängliga användarordlistorna.  
Markera användarordlistorna som du vill använda för rättstavningskontroll och avstavning.  
Ny  
Om du klickar på den här kommandoknappen kommer du till dialogrutan Skapa användarordlista där du gör inställningarna för den nya användarordlistan.  
Skapa användarordlista  
I området Ordlista kan du ge en ny användarordlista eller undantagsordlista ett namn och definiera språket.  
Namn  
Här anger du namnet på den nya användarordlistan.  
Filnamnstillägget "*.DIC" bifogas automatiskt.  
Språk  
Genom att välja ett visst språk begränsar du användningen av användarordlistan.  
Om du väljer Alla används användarordlistan oberoende av det aktuella språket.  
Undantag (-)  
Om du vill undvika vissa ord i dina dokument, markerar du den här rutan.  
I användarordlistan som definieras på det här sättet kan du lägga till alla ord som ska undvikas.  
Vid rättstavningskontrollen får du information om att ordet ska undvikas om den här undantagsanvändarordlistan är aktiverad.  
Redigera  
Om du klickar på den här kommandoknappen visas dialogrutan Redigera användarordlista där du kan utöka din användarordlista eller redigera poster som redan finns.  
I den här dialogrutan har du möjlighet att mata in nya ord eller redigera existerande poster.  
Om du redigerar en undantagsordlista finns det även möjlighet att definiera ett undantag för ett ord i dialogrutan.  
Vid en rättstavningskontroll kommer sedan det här undantaget upp som förslag.  
När du redigerar en ordlista kontrolleras vilken status filen har.  
Om den t.ex. är skrivskyddad går den inte att ändra.  
Kommandoknapparna Nytt och Radera är då deaktiverade.  
I så fall måste du första ändra filens status.  
I en nätverksinstallation av %PRODUCTNAME kan några användarordlistor ligga på servern i katalogen {installpath} / share / wordbook {installpath }\share\wordbook.  
De har installerats av systemadministratören, är skrivskyddade och innehåller t.ex. de ord som används specifikt på ditt företag.  
Dina egna användarordlistor ligger däremot i katalogen {installpath} / user / wordbook {installpath }\user\wordbook och går att redigera.  
Bok  
Här väljer du ut boken som du vill redigera.  
I ignorera-listan med namnet IgnoreAllList (Alla), som bara administreras för den aktuella rättstavningskontrollen i RAM-minnet, läggs alla ord till som du har markerat med Ignorera vid rättstavningskontrollen.  
Dessutom läggs en del av dina användardata (t.ex. namn, företag, gatuadress) till i listan vid programstarten.  
Det går inte att radera IgnoreAllList (Alla).  
Det går inte att välja bort posten IgnoreAllList och den kan inte raderas.  
Det går bara att radera orden som har lagts till som innehåll.  
Detta sker automatiskt varje gång du avslutar %PRODUCTNAME.  
Språk  
Här tilldelar du den aktuella användarordlistan ett nytt språk.  
Ord  
Här kan du mata in ett nytt ord som ska läggas till i ordlistan.  
I listrutan visas innehållet i den aktuella användarordlistan.  
Om du markerar ett ord från den här listan visas det i textfältet.  
Om du matar in ett ord med ett likhetstecken efter det, t.ex. AutoComplete=, varken avstavas det här ordet automatiskt eller föreslås för avstavning.  
Om du i stället matar in tecknet enligt mönstret Auto=Complete avstavas ordet bara på det här stället resp. föreslås för avstavning.  
Förslag  
Det här inmatningsfältet är bara tillgängligt om du redigerar en undantagsordlista.  
Fältet lägger till det alternativa förslaget till ordet i textfältet "Ord".  
Du gör så här med de båda textfälten för redigering av en undantagsordlista: anta att du alltid skriver "e-mail" som det är skrivet här.  
Vid korrigeringen vill du ha "email" som alternativ.  
Skriv e-mail i textfältet Ord och email i fältet Förslag.  
Nytt  
Klicka på den här kommandoknappen om du vill lägga till ordet som står i textfältet Ord och vid undantagsordlistor även ordet som står i fältet Förslag till din aktuella användarordlista.  
Radera  
Klicka på kommandoknappen Radera om du vill ta bort det markerade ordet från den aktuella användarordlistan.  
Radera  
Om du klickar på Radera kan du radera det markerade ordet efter en säkerhetskontroll såvida det inte är skrivskyddat.  
Alternativ  
I det här området definierar du alternativen för rättstavningskontrollen och avstavningen.  
Redigera  
Om du vill ändra ett värde, markerar du posten och klickar på Redigera.  
En dialogruta visas där du anger det nya värdet.  
Kontrollera ord med stora bokstäver  
Markera den här rutan om ord som bara innehåller stora bokstäver ska kontrolleras.  
Kontrollera ord med siffror  
Markera den här rutan om ord som förutom bokstäver även innehåller siffror ska kontrolleras.  
Kontrollera stor och liten bokstav  
Markera den här rutan om även den korrekta användningen av stora bokstäver i början av ord ska kontrolleras vid rättstavningskontrollen.  
Kontrollera specialområden  
Markera den här rutan om även specialområden, som t.ex. texter i sidhuvuden och sidfötter, i textdokumenttabeller och i textramar, ska kontrolleras vid rättstavningskontrollen.  
Kontrollera alla språk  
Om du markerar här värderas en överensstämmelse mellan ett ord och något av de installerade språken som korrekt.  
Teckenattributet "Språk" gäller alltså inte.  
Automatisk kontroll  
Om den här funktionen är aktiv, är den automatiska rättstavningskontrollen aktiverad.  
Eventuella felstavade ord stryks under med en röd korrekturlinje i ditt dokument.  
Om markören befinner sig på ett ord med en sådan markering och du öppnar snabbmenyn, visas en lista med ändringsförslag.  
Om du väljer något av förslagen, ersätter detta det markerade ordet.  
Om samma skrivfel återkommer senare i dokumentet, korrigeras det automatiskt.  
De automatiska ersättningarna gäller bara tills du avslutar %PRODUCTNAME.  
Om du vill föra in ordparet i ersättningstabellen för AutoKorrigering väljer du menykommandot AutoKorrigering på snabbmenyn för den automatiska korrigeringen.  
Välj ett förslag på undermenyn.  
Ordet ersätts och samtidigt förs ordparet in i ersättningstabellen.  
Dölj felmarkering  
Markera den här rutan om du vill att de röda våglinjerna ska döljas som indikerar rättstavningsfel när automatisk kontroll är aktiverad.  
I det här läget kontrolleras stavningen "i bakgrunden" medan du skriver eller när en text laddas, men den tidskrävande markeringen av felstavade ord utgår.  
Om du senare avmarkerar fältet Dölj felmarkering visas de röda linjerna direkt.  
Gammal tysk rättstavning  
Markera den här rutan om du bara vill använda den gamla tyska rättstavningen.  
Om rutan inte är markerad, använder %PRODUCTNAME de nya stavningsreglerna för rättstavningskontroll och avstavning.  
Minimal ordlängd för avstavning  
Ett ord avstavas aldrig automatiskt om det innehåller färre tecken än vad du ställer in här.  
Ange den minimala ordlängden i det här rotationsfältet eller antalet tecken före eller efter brytning.  
Tecken före radbrytning  
Den angivna siffran definierar hur många tecken som minst måste återstå av ett avstavat ord i slutet av raden.  
Tecken efter radbrytning  
Antalet bokstäver per stavelse som är angivet i textfältet definierar hur många bokstäver av ett avstavat ord som minst måste stå i början av nästa rad.  
Automatisk avstavning  
Om den här rutan är markerad blir du aldrig ombedd att göra ett manuellt avstavningsförslag.  
Om rutan inte är markerad öppnas en dialogruta där du kan avstava ord vars avstavning inte är känd.  
Avstava specialområden  
Om den här rutan är markerad avstavas ord även i fotnoter, sidhuvuden och sidfötter.  
Redigera moduler  
Här redigerar du modulerna.  
Alternativ  
I det här området väljer du ett språk och de moduler, som är aktiverade för det här språket, för rättstavning, avstavning och synonymordlista och du kan ordna modulerna efter prioritet.  
Välj först språk.  
Markera sedan alla moduler, som ska vara aktiverade för det här språket, under överskrifterna Rättstavning, Avstavning och Synonymordlista.  
När mer än en underordnad modul är tillgänglig för ett område bearbetas de underordnade modulerna för rättstavning och synonymordlista i den ordning som de står i listrutan.  
Du kan ändra ordningen med kommandoknapparna Prio + och Prio -.  
Vid avstavningen kan bara en enda underordnad modul vara aktiverad.  
Språk  
Här väljer du språk.  
Det står en bock framför en språkpost om det finns en rättstavningsmodul för det här språket.  
För alla andra språkurvalsfält i %PRODUCTNAME gäller följande:  
Det står en bock framför en språkpost om rättstavningskontrollen har aktiverats för det här språket.  
Prio +  
Om du klickar här höjer du prioriteten för modulen som är markerad i listrutan med ett steg.  
Prio -  
Om du klickar här minskar du prioriteten för modulen som är markerad i listrutan med ett steg.  
Tillbaka  
Klicka här om du vill ångra de aktuella ändringarna i listrutan.  
Färger  
Här kan du välja en färg från en färgtabell, ändra den och definiera nya färger.  
Färgtabell  
Namn  
Här kan du mata in ett nytt namn.  
Med Ändra ändras namnet på den aktuella färgen, med Lägg till definieras en ny färg.  
Färg  
Här väljer du en färg.  
Färgmodell  
Färgmodell  
Här väljer du färgmodell:  
Röd-Grön-Blå (RGB) eller Cyan-Magenta-Yellow-Black (CMYK).  
Bredvid dem kan du i ett rotationsfält definiera värdet för respektive färg från 0 till 255.  
R  
Välj andelen rött.  
G  
Välj andelen grönt.  
B  
Välj andelen blått.  
Bredvid dem kan du i ett rotationsfält definiera värdet för respektive färg från 0 till 255.  
C  
Välj andelen cyan.  
M  
Välj andelen magenta.  
Y  
Välj andelen gult (yellow).  
K  
Välj andelen svart (black).  
Lägg till  
Med den här kommandoknappen lägger du till en ny färg.  
Ändra  
Med den här kommandoknappen ändrar du den aktuella färgen.  
Någon säkerhetskontroll sker inte, färgen skrivs över.  
Redigera...  
Ladda färgtabell  
Med den här ikonen kommer du till dialogrutan Öppna där du kan öppna en färgtabell.  
Spara färgtabell  
Med den här ikonen öppnar du dialogrutan Spara som, där du kan spara den aktuella färgtabellen med ett eget namn.  
Om du inte väljer det här kommandot, sparas den aktuella färgtabellen automatiskt som standard och laddas automatiskt igen när du startar %PRODUCTNAME nästa gång.  
Ikonerna Ladda färgtabell och Spara färgtabell visas bara om du öppnar fliken Färger via kommandot Format - Yta....  
Färg  
Här kan du definiera en egen färg i en tvådimensionell tonad grafik och / eller numeriskt.  
Den nya färgen visas i det undre förhandsvisningsfältet på sidan Färger när du har stängt den här dialogrutan med OK.  
Där kan du bestämma om du vill lägga till färgen i den aktuella färgpaletten som en helt ny färg eller om den nya färgen ska ersätta färgen som visas i det övre förhandsvisningsfältet.  
Färgfönster  
I de båda stora färgfönstren väljer Du en ny färg genom att klicka på den med musen.  
Du kan välja färg både från det vänstra och det högra färgfönstret.  
I det högra färgfönstret visas hela färgspektrumet från vänster till höger.  
I den över delen av fönstret är färgerna helt mättade och i den undre är de omättade.  
I det vänstra färgfönstret visas ett urval av färger som visar ett stegvis uppdelat spektrum mellan de fyra färgerna i hörnen av fönstret.  
Du ändrar färgerna i de fyra hörnen på följande sätt:  
Klicka i hörnfältet vars färg du vill ändra.  
Du kan också definiera färgen genom att ange värden i de numeriska inmatningsfälten.  
Överför färgen som du har valt till höger till det lilla fältet som är markerat i det vänstra färgfönstret genom att klicka på kommandoknappen <- -.  
Färggradienten i det vänstra färgfönstret anpassas direkt i färgton, mättnad och ljusstyrka.  
<- -  
Överför den färg som du har valt till höger till hörnfältet som är markerat i det vänstra färgfönstret genom att klicka på kommandoknappen <--.  
-->  
Placerar den lilla urvalsmarkören i det högra fönstret på den färg som motsvarar den markerade färgen i det vänstra fönstret och uppdaterar värdena i de numeriska inmatningsfälten.  
Cyanblått  
Här väljer Du färgvärdet cyan i CMYK-färgmodellen.  
Magenta  
Här väljer du färgvärdet Magenta i CMYK-färgmodellen.  
Gult  
Här väljer du färgvärdet gult (yellow) i CMYK-färgmodellen.  
Key  
Key (svart) i CMYK-färgmodellen.  
Rött  
Här väljer du färgvärdet rött i RGB-färgmodellen.  
Grönt  
Här väljer du färgvärdet grönt i RGB-färgmodellen.  
Blått  
Här väljer du färgvärdet blått i RGB-färgmodellen.  
Färg  
Här väljer du färgton (hue) i HSB-färgmodellen.  
Mättnad  
Här väljer du mättnad (saturation) i HSB-färgmodellen.  
Ljusstyrka  
Här väljer du ljusstyrka (brightness) i HSB-färgmodellen.  
I det vänstra förhandsvisningsfältet visas originalfärgen från den överordnade sidan Färger.  
I det högra förhandsvisningsfältet visas alltid det aktuella resultatet av ditt arbete i den här dialogrutan.  
Allmänt  
Här gör du allmänna inställningar för %PRODUCTNAME.  
Tvåsiffriga årtal  
Här väljer du intervallet som ska gälla vid inmatning av tvåsiffriga årtal.  
Årtalen i datumangivelser angavs tidigare för det mesta med två siffror.  
Internt hanterar %PRODUCTNAME årtal med fyra tecken, vilket innebär att programmet korrekt kan beräkna tiden mellan den 1 / 1 99 till den 1 / 1 01 till två år.  
Här kan du ställa in till vilket år ett tvåsiffrigt årtal ska adderas till 2000.  
Det förvalda värdet är det gränsvärde som är inställt i operativsystemet, t.ex. "30".  
Det innebär att om du anger 1 / 1 30 eller ett senare datum, behandlas det internt som 1 / 1 1930 eller senare.  
Det innebär att den 1 / 1 20 tolkas som den 1 / 1 2020.  
Help Agent  
I det här området bestämmer du hur Help Agent ska fungera.  
Aktivera  
Om den här rutan är markerad visas Help Agent automatiskt i utvalda situationer.  
Visningstid  
Välj här hur länge Help Agent ska visas innan den stängs automatiskt.  
Återställ Help Agent  
Om du inte har öppnat Help Agent i en viss situation tre gånger efter varandra, utan stängt den eller låtit den stängas automatiskt, visas Help Agent aldrig mer i den här situationen.  
Situationen tas bort från den interna listan.  
Om du klickar här återställs listan med situationerna då Help Agent visas till grundinställningen.  
Öppna / spara-dialogrutor  
Använd %PRODUCTNAME -dialogrutor  
Om du markerar den här rutan används %PRODUCTNAME -dialogrutorna när dokument ska öppnas och sparas, i annat fall operativsystemets dialogrutor.  
I %PRODUCTNAME -hjälpen beskrivs %PRODUCTNAME -dialogrutorna för att Öppna och Spara dokument.  
Dokumentstatus  
Utskrift sätter status "~Dokument ändrat"  
Om den här rutan är markerad gäller utskrift av dokument som ändring.  
Det innebär att du blir tillfrågad om ändringarna ska sparas när du har sparat och skrivit ut ett dokument och stänger det direkt efter det.  
I så fall registreras utskriftsdatum som ändring i dokumentegenskaperna.  
Teckensnittsersättning  
Här kan du påverka de teckensnitt som ditt system ställer till förfogande för %PRODUCTNAME.  
Om ett teckensnitt inte går bra att läsa på ditt system väljer du ett annat teckensnitt och markerar fälten "Alltid" och "Bildskärm ".  
Även vid laddning av externa dokument (t.ex. HTML-dokument) kan ersättningen av teckensnitt vara till hjälp.  
Om teckensnittet i den laddade filen inte finns på ditt system, avgör systemet vilket teckensnitt som ska användas i stället.  
Om du inte vill ha det kan du ersätta det.  
Ersättningen av teckensnitt ändrar inte dokumenten utan gäller bara den datormiljö som används.  
Använd ersättningstabell  
Med den här rutan definierar du om ersättningstabellen som du har skapat ska användas.  
Ersättningstabell  
När du har valt och övertagit ett teckensnittspar, visas både originalteckensnittet och ersättningsteckensnittet här.  
Ändringarna gäller dokument, dialogrutor och så vidare.  
Alltid  
Markera den här rutan om du vill att originalteckensnittet ska ersättas även om det finns på ditt system.  
Ett dokument som ursprungligen sparades med Times New Roman, visas med det nya teckensnittet även om Times New Roman är installerat i ditt system.  
Om Alltid inte är markerat, ersätts bara de teckensnitt som inte finns i ditt system.  
Om exempelvis teckensnittet Times New Roman finns i ditt system, och Alltid inte är markerat, ersätts aldrig det här teckensnittet.  
Bildskärm  
Om den här rutan är markerad, gäller ersättningen av teckensnitt bara bildskärmen och inte utskrift.  
Har du en Postscript-skrivare och använder ett system som även har TrueType-teckensnitt?  
Om du vill att utskrifter å ena sidan alltid ska göras med Postscript-teckensnitt, men visningen på bildskärmen å andra sidan alltid med TrueType-teckensnitt, gör du som i följande exempel:  
Alltid  
Bildskärm  
Teckensnitt  
Ersätt med  
aktivera  
deaktivera  
Arial  
Helvetica  
aktivera  
deaktivera  
Times New Roman  
Times  
aktivera  
deaktivera  
Courier New  
Courier  
Vid HTML-filer kan du förbättra ersättningen av teckensnitt om du markerar rutan Ignorera teckensnittsinställningar i dialogrutan som öppnas med menykommandot Verktyg - Alternativ - Ladda / spara - HTML-kompatibilitet.  
Teckensnitt  
Använd det här kombinationsfältet till att ange eller välja ut teckensnittet som ska bytas ut.  
Ersätt med  
I det här kombinationsfältet anger du ersättningsteckensnittet.  
Du kan mata in det direkt eller välja ut det i listan.  
Överta  
Klicka här om du vill överta det aktuella teckensnittsparet till listrutan.  
Överta  
Radera  
Klicka här om du vill radera det markerade teckensnittsparet från listan.  
Radera  
Vy  
Här finns fler inställningsmöjligheter för vyn.  
Visning  
Utseende  
I det här kombinationsfältet kan du göra %PRODUCTNAME mer likt andra operativsystem.  
Standard  
Det här är standardinställningen och den visar fönster, kryssrutor o.s.v. enligt Sun Microsystems förinställningar.  
Macintosh  
Om du vill att %PRODUCTNAME ska påminna om en Apple-Macintosh när du arbetar, väljer du den här posten.  
XWindows  
Om du väljer den här posten ser %PRODUCTNAME som XWindows.  
OS / 2  
Välj den här posten om du vill att %PRODUCTNAME ska se ut som OS / 2.  
Skalning  
I det här rotationsfältet ställer du in en procentuell storleksförändring för bildskärmsvisningen av teckenstorleken.  
De ändringar som du gör här påverkar storleken på all text på skärmen (t.ex. text i dialogrutor, ikonetiketter).  
Inställningen Skalning har inte något med den faktiska teckenstorleken i dina texter att göra.  
Det är bara fråga om en förstorad visning på bildskärmen.  
Återställ  
Här kan du bestämma vilken redigeringsvy för dokument och fönster som ska återställas när du startar %PRODUCTNAME på nytt.  
Redigeringsvy  
Här definierar du om den senast använda dokumentvyn, som du valde i %PRODUCTNAME, ska återställas.  
De egenskaper som gällde då du senast sparade dokumentet återställs.  
För textdokument gäller det bl.a. markörens läge, för tabelldokument den tabell och fönsteruppdelning som visas, för presentationsdokument det valda sidläget eller bakgrundsläget.  
Öppnade fönster  
Här definierar du om de fönster som är öppna när programmet avslutas ska återställas när %PRODUCTNAME startas igen.  
Jämna ut bildskärmsteckensnitt (antialiasing)  
Om du markerar den här rutan jämnas bildskärmsteckensnitten ut.  
I rotationsfältet ställer du in från och med vilken storlek i pixel teckensnitten ska jämnas ut.  
Meny följer muspekaren  
Om den här rutan är markerad följer markeringen av en meny resp. undermeny med när du flyttar muspekaren.  
Registerkort på en rad  
Om du markerar den här rutan visas registerkort i dialogrutor med många registerkort på en rad.  
Registerflikar i färg  
Markera den här rutan om du vill ha registerflikar i färg.  
Förhandsvisning i teckensnittslistor  
Om du markerar den här rutan visas namnen på teckensnitten formaterade med respektive teckensnitt, t.ex. i fältet Teckensnitt på objektlisten.  
Inaktiva menyposter  
Om du markerar den här rutan visas alla inaktiva menyposter i grått.  
Om rutan inte är markerad döljs alla menykommandon som inte är tillgängliga.  
Teckensnittshistorik  
De visas i kombinationsfältet Teckensnittsnamn på objektlisten.  
Upp till 5 teckensnitt visas och det senast använda teckensnittet infogas alltid överst i listan.  
Stora ikoner  
Om den här rutan är markerad förstoras ikonerna på symbollisterna.  
Flata ikoner  
Markera den här rutan om du vill att ikonerna på symbollisterna ska vara flata.  
Visa ikoner på menyer  
Om den här rutan är markerad visas de tillhörande ikonerna framför respektive menypost.  
3D-visning  
Använd OpenGL  
Om den här rutan är aktiv visas 3D-grafik från %PRODUCTNAME Draw och %PRODUCTNAME Impress med hjälp av den hårdvara som stöder OpenGL i systemet.  
Om ditt system inte innehåller någon hårdvara som stöder OpenGL, ignoreras inställningen i den här rutan.  
Om du avmarkerar rutan görs 3D-visningen alltid per program.  
Optimerad utmatning  
Om det här fältet är markerat får du en optimerad OpenGL-utmatning.  
Om "Optimerad utmatning" är aktiverat överförs all geometridata samtidigt i en matris till grafikdrivrutinen.  
Men det är inte alla grafikdrivrutiner som stödjer denna OpenGL-funktion på rätt sätt.  
Därför kan du avmarkera "Optimerad utmatning" om det uppstår fel i samband med 3D-visning.  
Det innebär att all geometridata överförs som enskilda punkter efter varandra.  
Använd ditrering  
Använd det här alternativet om Du vill att få färger ska visas som om det fanns fler färger.  
Ditreringsfunktionen utnyttjar det faktum att det mänskliga ögat uppfattar två färgpunkter (pixlar) som ligger alldeles intill varandra, som en blandning av båda.  
En schackbrädesliknande blandning av svarta och vita punkter gör att det mänskliga ögat uppfattar ytan som grå.  
Det här alternativet aktiveras som standard.  
De används för att ditrera framställningar med färre färger.  
Eftersom många bitar av färginformationen faller bort utan ditrering är effekten av en sådan gradering mycket tydlig.  
Kvaliteten blir sämre ju färre färger som används.  
Full visning vid interaktion  
Istället ser du en full visning av 3D-objektet.  
Standardinställningen är att alternativet är avmarkerat.  
Musplacering  
Här väljer du om och hur muspekaren placeras i en dialogruta när den öppnas.  
Musknapp i mitten  
Här väljer du hur musknappen i mitten ska fungera.  
Automatisk rullning - om du håller ner musknappen i mitten och drar i ett dokument flyttas vyn.  
Infoga urklipp - om du klickar med musknappen i mitten infogas innehållet i "Selection Clipboards" urklippet vid markörens position.  
Urklipp  
Selection Clipboard  
Definiera innehåll  
Redigera - Kopiera Ctrl+C.  
Markera text, tabell, objekt.  
Klistra in innehåll  
Redigera - Klistra in Ctrl+V infogar vid textmarkörens position.  
Klick med musknappen i mitten klistrar in vid muspekarens position.  
Vid dokumentbyte  
Ingen påverkan av innehållet i urklippet.  
Den markering som är synlig senast är innehållet i Selection Clipboards.  
Skriv ut  
Här hittar du inställningsmöjligheter för utskrift.  
Reducera utskriftsdata  
I det här området definierar du att färre data överförs till skrivaren.  
När utskriftsdata reduceras skriver skrivaren ut snabbare, även laserskrivare kan skriva ut med mindre minne och mindre utskriftsfiler skapas.  
Nackdelen är att utskriftskvaliteten blir sämre.  
Inställningar för  
Välj här om de följande inställningarna i det här området ska gälla för direkt utskrift på skrivaren eller för utskrift till en fil.  
Reducera transparens  
Om du markerar den här rutan skrivs transparenta objekt ut som normala, icke-transparenta objekt, beroende på vad du väljer i de båda följande alternativfälten.  
Transparens kan för närvarande inte matas ut på någon skrivare.  
Områdena i ett dokument där det finns transparens måste därför alltid beräknas som bitmap och skickas till skrivaren.  
Beroende på bitmapstorlek och utskriftsupplösning kan det uppstå väldigt mycket data på det här sättet.  
Automatiskt  
Med det här alternativet skrivs bara transparensen ut när den transparenta ytan täcker mindre än en fjärdedel av hela sidan.  
Ingen transparens  
Med det här alternativet skrivs transparens aldrig ut.  
Reducera bitmaps  
Om du markerar den här rutan skrivs bitmaps ut i reducerad kvalitet.  
Upplösningen kan bara minskas, inte höjas.  
Hög / Normal utskriftskvalitet  
Hög utskriftskvalitet motsvarar en upplösning på 300 dpi.  
Normal utskriftskvalitet motsvarar en upplösning på 200 dpi.  
Upplösning  
Med det här alternativet bestämmer du själv den maximala utskriftskvaliteten i dpi.  
Upplösningen kan bara minskas, inte höjas.  
Inkludera transparenta objekt  
Om den här rutan är markerad gäller reduceringen av utskriftskvalitet för bitmaps även för transparenta områden i objekt.  
Reducera färggradienter  
Om den här rutan är markerad skrivs färggradienter ut i reducerad kvalitet.  
Färggradientränder  
Här väljer du det maximala antalet färggradientränder för utskrift.  
Mellanfärg  
Med det här alternativet skrivs färggradienter bara ut i en mellanfärg.  
Omvandla färger till gråskalor  
Om den här rutan är markerad skrivs alla färger bara ut som gråskalor.  
Skrivarvarningar  
Här ställer du in vilka varningar som ska visas innan utskriften påbörjas.  
Pappersstorlek  
Markera den här rutan om du behöver en speciell pappersstorlek när du skriver ut det aktuella dokumentet.  
Om den aktuella skrivaren inte har den pappersstorlek som används i dokumentet får du ett felmeddelande.  
Pappersorientering  
Markera den här rutan om du behöver en speciell pappersorientering när du skriver ut det aktuella dokumentet.  
Om den aktuella skrivaren inte har den pappersorientering som används i dokumentet får du ett felmeddelande.  
Transparens  
Markera den här rutan om du alltid vill varnas när ett dokument innehåller transparenta objekt.  
Om du skriver ut ett sådant dokument visas en dialogruta, där du kan välja om transparensen ska skrivas ut i det här utskriftsjobbet eller inte.  
Här öppnar du en dialogruta där du kan söka efter program.  
Hjälpprogram  
Här kan du ange vilket program som ska utföra vilken tjänst.  
Skicka dokument som e-post med  
I det här området definierar du med vilket program ett dokument skickas som e-post när du väljer kommandot under Arkiv - Skicka.  
Även när du klickar på en mailto:-URL i ett dokument startas det program som har valts här.  
Standardprogram för e-post  
Markera den här rutan om det program som är registrerat som standardprogram för e-post i ditt system ska startas när du vill skicka e-post från %PRODUCTNAME.  
Om du arbetar med Netscape 4.7x som e-postprogram i Unix, är det bäst att använda skriptet nswrapper som ligger i katalogen {installpath} / program.  
Om Netscape 4.7x finns i sökvägen behöver du inte ändra skriptet.  
Andra  
Här väljer du ett program som e-postprogram.  
Profiler  
Välj en profil.  
Profilen definierar på vilket sätt parametrar ska överföras till programmet.  
Program  
Mata in programmets sökväg och namn eller klicka på... och välj ut det i dialogrutan som öppnas.  
Utför länkar med  
Här väljer du programmet som används för en tjänst när den startas via en länk i ett dokument.  
HTTP  
Välj program för protokollet HTTP.  
HTTPS  
Välj program för protokollet HTTPS.  
FTP  
Välj program för protokollet FTP.  
MAILTO  
Välj program för protokollet SMTP.  
Filhanterare  
Här väljer du filhanterare.  
Den startas om en fil öppnas från %PRODUCTNAME som %PRODUCTNAME inte kan öppna själv, eftersom filtypen inte är känd i %PRODUCTNAME.  
Program  
Mata in programmets namn och sökväg eller klicka på... och välj det i dialogrutan som öppnas.  
Arbetsminne  
Här gör du bl.a. förinställningarna för grafikcachen, bestämmer hur många steg som går att ångra samt om du vill använda snabbstart av %PRODUCTNAME.  
Ångra  
Här ser du hur många steg som du maximalt kan ångra.  
Antal steg  
I det här rotationsfältet väljer du antalet steg som ska gå att ändra.  
Grafikcache  
Grafikcachen sparar den grafik som ett dokument innehåller i arbetsminnet på din dator.  
Du kan visa samma grafik direkt, t.ex. när du har rullat i dokumentet, utan att t.ex. skalning, sektion, filter o.s.v. måste beräknas om igen.  
Använd för %PRODUCTNAME (MB)  
Välj den totala cachestorleken för all grafik.  
Minne per objekt (MB)  
Objekt som är större än vad du väljer här lagras inte i cachen.  
Ta bort från minnet efter (hh:mm)  
Här väljer du hur länge varje grafikobjekt finns kvar i cachen i timmar och minuter.  
Cache för infogade objekt  
Antal objekt  
Välj här det maximala antalet OLE-objekt som lagras i cachen.  
Snabbstart av %PRODUCTNAME  
Ladda %PRODUCTNAME vid systemstart  
Markera den här rutan om %PRODUCTNAME ska förberedas för snabbstart när systemet startar.  
Om snabbstarten är aktiverad laddas delar av %PRODUCTNAME i minnet redan när systemet startar.  
På aktivitetsfältet finns en ikon vars snabbmeny bl.a. innehåller kommandon som du kan öppna %PRODUCTNAME -dokument med.  
Alternativ Ladda / spara  
Här gör du allmänna inställningar som gäller när du laddar / sparar.  
Proxy  
Här gör du inställningar för proxyservrar.  
Proxyservrar används för åtkomst till Internet via ett mellanliggande nätverk och kan antingen konfigureras automatiskt eller manuellt.  
Inställningar  
I det här området gör du inställningarna som du behöver för att kommunicera med Internet via en proxyserver.  
Proxyserver  
I den här listrutan väljer du typ av proxydefinition.  
Ingen  
Välj det här alternativet om åtkomsten till Internet sker utan proxyserver.  
Detta är fallet när du skapar en förbindelse direkt från arbetsdatorn till en Internet-leverantör som inte använder någon proxyserver.  
Manuellt  
Välj den här posten om du själv måste ange de nödvändiga och / eller önskade proxyservrarna.  
Du kan specificera proxyservrarna i de textfält som följer.  
Proxyservrarna måste eventuellt anropas på olika sätt, beroende på Internet-tjänst.  
Fråga systemadministratören vilka data du ska ange här.  
I textfälten i den här dialogrutan anger du servernamn utan protokollbeteckningen: www.sun.com är t.ex. rätt, men inte http: / /www.sun.com.  
Http proxy  
I det här textfältet anger du namnet på proxyservern för HTTP (webbsidor).  
Porten anger du i det högra fältet.  
Ftp proxy  
I det här textfältet anger du namnet på proxyservern för FTP.  
Porten anger du i det högra fältet.  
Socks proxy  
I det här textfältet anger du namnet på proxyservern för Socks.  
Porten anger du i det högra fältet.  
Ingen proxy för:  
Ange här namnen på de servrar där inga proxyservrar ska användas.  
Det är t.ex. de servrar som ska anropas i det egna lokala nätverket och servrar vars kapacitet skulle minska om de mellanlagras via en proxy (t.ex. video - och audio-direktförbindelser, webbkameror).  
Avgränsa namnen med semikolon (;).  
Du kan alltså t.ex. ange "*.sun.se" (utan citattecken) om alla värddatorer i domänen sun.se ska anropas utan proxy, eller "www.lifevideo.* "för att anropa alla www.lifevideo-värddatorer utan proxy i hela världen (detta är ett fiktivt exempel).  
Port  
I textfälten anger du porten för respektive proxyserver som står bredvid.  
Det högsta värdet som kan anges för en port är 65535.  
DNS-server  
Här ställer du in DNS (Domain Name System).  
DNS-namnservern används till att omvandla det fullständiga namnet på den dator, som du anger i en URL (t.ex. www.sun.se), till dess 32 bitars IP-adress.  
32-bit-talen i IP-adresser visas för översiktlighetens skull i fyra decimaltal som är förbundna med punkter.  
Varje decimaltal ligger mellan 0 och 255 och representerar de första, andra, tredje och sista 8 bitarna av de totala 32 bitarna.  
Automatiskt  
Automatisk överföring av DNS från systeminställningarna.  
Den här inställningen rekommenderas.  
När du går in på Internet via anslutningar med olika leverantörer kan du t.ex. automatiskt använda den namnserver som leverantören rekommenderar (vars IP-adress du t.ex. har angett i DFÜ-nätverksdialogrutan).  
Manuellt  
Manuell inmatning av DNS.  
Ange IP-adressen för DNS-servern i textfältet med det vanliga skrivsättet för IP-adresser.  
Sökning  
Här definierar du hur %PRODUCTNAME ska använda sökmotorerna på Internet.  
Sök i  
I det här området anger du dina alternativ.  
I de följande exemplen används www.altavista.com i den version som var giltig när den här texten skrevs.  
När du läser den här texten kan Altavista ha ändrats - anpassa dig i så fall efter det när du använder exemplet. "AltaVista® is a registered trademark of AltaVista Company."  
Sökmotorer  
I den här listrutan visas sökmotorerna som redan är definierade.  
Om du markerar en av sökmotorerna, visas respektive konfiguration i text - och alternativfälten som finns bredvid.  
Namn  
I det här textfältet kan du föra in namnet på en sökmotor.  
Det är det namn som visas på undermenyn till ikonen Sök.  
Typ  
I det här alternativområdet väljer du ut för vilken typ av sökordskombinationer som konfigurationen i textfälten nedanför ska definieras eller visas.  
Du kan välja mellan Och, Eller och Exakt.  
Du måste alltid definiera alla tre alternativen fullständigt och klicka på kommandoknappen Ändra efter varje ändring.  
Prefix  
I det här textfältet skrivs eller visas webbadressen och den första delen av sökkommandot för en sökmotor.  
Om du söker med av de HTML-baserade Internet-sökmotorerna, t.ex. efter "%PRODUCTNAME" med Altavista, visas den kompletta URL:en för den här sökningen i URL-inmatingsfältet i din webbläsare.  
Du får följande URL för det här exemplet:  
http: / /www.altavista.com / cgi-bin / query?q= %PRODUCTNAME &kl=XX&pg=q&Translate=on  
I fältet Prefix kopierar du allt som står framför söktexten, följande i det här exemplet:  
http: / /www.altavista.com / cgi-bin / query?q=  
Detta är den första delen av sökfrågan.  
Om du har angett flera ord som är åtskilda med mellanslag, infogas det tecken som finns i fältet Skiljetecken för att koppla ihop orden.  
Suffix  
Sökorden placeras mellan prefixet och suffixet.  
Suffixet anger den kommandosekvens som skickas i slutet av ett sökkommando.  
I det här exemplet är det följande:  
&kl=XX&pg=q&Translate=on  
Skiljetecken  
Om du anger flera ord i en sökning, skiljs de åt med tecknen som är angivna i det här textfältet.  
De flesta sökmotorer kräver här ett plustecken (+).  
Så här tar du reda på vilka prefix, skiljetecken och suffix som du måste ange när du definierar en ny sökmotor.  
Gå till sökmotorn och gör en sökning med minst två ord.  
Kopiera webbadressen från fältet URL på funktionslisten och klistra in den i ett tomt dokument.  
Ändra villkoret för sökningen i sökmotorn, om det finns möjlighet att välja.  
Kopiera innehållet i fältet URL en gång till.  
Jämför webbadresserna med exempeladresserna, som Du kan kopiera från fälten i den här dialogrutan.  
Du bör sedan kunna urskilja prefix, suffix och skiljetecken för respektive villkor.  
Skrivstil  
I den här listrutan väljer du hur %PRODUCTNAME ska hantera stor och liten bokstav i sökorden.  
Posterna är Liten, Stor och Ingen.  
Beroende på vilken post du väljer görs sökorden om till gemener, versaler eller inte alls.  
Många sökmotorer behandlar sökningar olika beroende på hur de är skrivna.  
Om du använder Altavista och skriver orden med små bokstäver, hittas alla ord oavsett om de är skrivna med stora eller små bokstäver.  
Men om sökordet däremot är skrivet med en eller flera versaler någonstans i ordet, hittas bara de ord som är skrivna exakt likadant.  
I vårt exempel med Altavista är det alltså bäst att inte omvandla skrivsättet (d.v.s. att välja Ingen).  
Nytt  
Med den här kommandoknappen lägger du till en ny sökmotor.  
Med Nytt raderar du alla poster som "Namn", "Suffix" och så vidare.  
Du måste alltså ange alla nödvändiga uppgifter för den nya sökmotorn från början.  
När du har övertagit uppgifterna med Lägg till visas den nya sökmotorn i listan över sökmotorer i området Sök i.  
Du kan börja använda den nya sökmotorn direkt.  
Lägg till  
Genom att klicka på den här kommandoknappen lägger du till en ny konfiguration i listan med konfigurationer.  
Ändra  
Om du har ändrat en konfiguration som redan är definierad, övertar du ändringarna med den här knappen.  
Radera  
Om du klickar på den här kommandoknappen, raderas den markerade sökmotorn direkt utan att du behöver bekräfta detta innan.  
Alternativ Internet  
Här gör du inställningar för Internet.  
Säkerhet  
Här definierar du om %PRODUCTNAME Basic-skript ska utföras.  
Om du begränsar listan med tillförlitliga URL:er eller väljer Kör makro - aldrig, visas eventuellt ett felmeddelande om att "rättigheter saknas" när du försöker köra ett skript, t.ex. när du försöker köra en AutoPilot eller ladda en mall.  
Standarden för tillförlitliga URL:er kan du återställa efter en eventuell ändring genom att klicka på kommandoknappen Standard.  
%PRODUCTNAME Basic-skript  
%PRODUCTNAME Basic-skript  
Här väljer du hur %PRODUCTNAME Basic-skript ska behandlas.  
Enligt sökvägslista  
Om du väljer det här alternativet, så utförs bara sådana %PRODUCTNAME Basic-skript som kommer från de URL:er som finns med i listrutan.  
Alltid  
Om du väljer det här alternativet, så utförs alla %PRODUCTNAME Basic-skript, oavsett ursprung.  
Aldrig  
Om du väljer det här alternativet, så utförs inte något %PRODUCTNAME Basic-skript alls, oavsett ursprung.  
Fråga vid andra dokumentkällor  
Om ett dokument, som du öppnar från en källa som inte finns med på listan, innehåller ett makro, blir du ombedd att bekräfta att makrot ska köras innan det körs.  
Om den här rutan inte är markerad körs makrot utan säkerhetsfråga.  
Visa varning innan makro körs  
Markera den här rutan om du vill bli varnad när ett makro körs.  
I en dialogruta tillfrågas du om %PRODUCTNAME Basic-makrona ska köras.  
Detta gäller också om ett dokument, som innehåller makroanrop i formler, laddas.  
Sökvägslista  
De tillförlitliga URL:erna visas i listrutan.  
Du kan markera och radera poster, eller återställa alla poster till standard.  
URL  
Innebörd  
$(workdirurl)  
Din arbetskatalog (se Verktyg - Alternativ - %PRODUCTNAME - Sökvägar).  
$(userurl)  
Vid en fristående installation är det $(insturl) / user.  
Vid en nätverksinstallation är det user-mappen under mappen till din användarinstallation.  
$(insturl)  
Vid en fristående installation är det {installpath} om du inte har ändrat det vid installationen.  
Vid en nätverksinstallation ligger installationskatalogen för det mesta på servern (se installationshandboken).  
Ny sökväg  
I textfältet skriver du en ny URL som du vill lägga till på listan med tillförlitliga URL:er.  
Du kan även använda jokertecken vid inmatningen, som t.ex. i *sun*.  
Klicka sedan på Lägg till.  
Om du anger en file: / / URL i filsystemet, är alltid alla underordnade kataloger inkluderade.  
Lägg till  
Klicka här om du vill lägga till en ny URL som du har angett i textfältet till listrutan.  
Frige  
Plug-ins  
Markera den här rutan om du vill att plug-ins ska kunna köras i dokument.  
Appletprogram  
Markera den här rutan om du vill att appletprogram ska kunna köras i dokument.  
Java  
I det här området väljer du hur Java-program ska behandlas.  
frige  
Om den här rutan är markerad kan Java-program köras.  
Extern Java-kod säkerhetskontrolleras automatiskt så länge rutan Säkerhetskontroller är aktiverad.  
Du får en varning om Java-kod upptäcks som vill komma åt din hårddisk.  
Säkerhetskontroller  
Om du deaktiverar den här rutan genomför Java inga säkerhetskontroller för extern kod (t.ex. appletprogram).  
Läs i varje fall följande information i hjälpen!  
Kod gäller som "extern" när den inte är tillgänglig via inställd ClassPath (se nedan).  
Appletprogram kan läsa och skriva på alla enheter om kontrollen inte är aktiverad!  
Eftersom JavaScript kan komma åt hela Java-miljön via LiveConnect-gränssnittet finns den här möjligheten även för JavaScript när kontrollen är avstängd.  
Stäng i varje fall av säkerhetskontrollerna om något av följande villkor är uppfyllt:  
Om du vet exakt vad appletprogrammet, Java-programmet eller JavaScript kommer att utföra,  
eller om du är inloggad som gästanvändare i Windows NT / 2000 eller Unix och du därför hindras att läsa och förstöra säkerhetsrelevanta data av operativsystemet.  
Nätåtkomst  
Här styr du Java-programs åtkomst till ditt nätverk.  
Du kan tillåta Obegränsad åtkomst, begränsa den till den aktuella Värddatorn eller förhindra den fullständigt med Ingen.  
ClassPath  
Med den här inställningen kan du lägga till fler Java-klasser eller Java-klassbibliotek för Java-miljön i %PRODUCTNAME.  
Enskilda sökvägar skiljs åt med;.  
Om kataloger finns med måste de avslutas med ett\ i slutet.  
Java-klasser som anropas via ClassPath säkerhetskontrolleras inte, i motsats till Java-klasserna som t.ex. anropas via en <APPLET>-tagg på en HTML-sida.  
...  
Med den här kommandoknappen kommer du till dialogrutan Välj sökvägar där du kan välja en ClassPath.  
HTML-kompatibilitet  
Här gör du inställningar för HTML-dokument.  
Teckenstorlekar  
Ställ in teckenstorlek i rotationsfälten Storlek 1 till Storlek 7 för visningen av taggarna <font size=1> till <font size=7>.  
Import  
I det här området gör du inställningar för import av HTML-dokument.  
Importera okända HTML-taggar som fält  
Aktivera den här rutan om du vill att taggar som %PRODUCTNAME inte känner igen ska importeras som fält.  
För en "normal" tagg i formen <Tag> skapas ett HTML_ON-fält med taggnamnets värde och för en avslutande tagg i formen < / Tag> skapas ett HTML_OFF-fält.  
Vid export till HTML omvandlas fälten till taggar igen.  
Ignorera teckensnittsinställningar  
Då används de teckensnitt som definierats i din HTML-sidformatmall.  
Export  
I det här området gör du inställningar för export av HTML-dokument.  
Vid export i HTML-format väljer du filtypen Webbsida i dialogrutan Spara som.  
Det finns mer information i beskrivningen av import - och exportfilter.  
Välj i kombinationsfältet för vilken standard eller webbläsare HTML-exporten från %PRODUCTNAME ska optimeras.  
HTML 3.2  
Om Du vill att HTML 3.2-specifika instruktioner ska beaktas vid export ska Du aktivera detta alternativ i listrutan.  
MS Internet Explorer 4.0  
Välj denna post i listrutan om Du vill att MS Internet Explorer 4.0-instruktioner ska beaktas vid export.  
Netscape Navigator 3.0  
Genom att aktivera denna post i listrutan beaktas bl a Netscape 3:s programtillägg multicol och Spacer vid export.  
Netscape Navigator 4.0  
Via denna post i listrutan aktiveras Netscape 4-programtillägg för export till HTML.  
Till skillnad från exportformatet %PRODUCTNAME Writer kan dock inte anfanger, små kapitäler, styckebakgrunder och kerninguppgifter exporteras.  
%PRODUCTNAME Writer  
Om Du vill att %PRODUCTNAME Writer-specifika instruktioner ska beaktas vid export ska Du aktivera detta alternativ i listrutan.  
StarBasic  
Om Du markerar detta fält så beaktas %PRODUCTNAME Basic-instruktioner vid export till HTML.  
Du måste aktivera det här alternativet innan du skapar ett %PRODUCTNAME Basic-skript, annars infogas det inte. %PRODUCTNAME Basic-skript måste stå i HTML-dokumentets huvud.  
När du har skapat makrot i %PRODUCTNAME Basic IDE visas det i källtexten i HTML-dokumentets huvud:  
Om makrot ska starta automatiskt när HTML-dokumentet öppnas, går du till dialogrutan Verktyg - Anpassa - Händelser och väljer "Dokument" uppe till höger i alternativrutan, "Öppna dokument "i händelselistan och väljer under Makron, ett dokument, dokumentets standardbibliotek, Modul1 och makrot.  
Klicka sedan på Tilldela.  
Visa varning  
Om den här rutan är markerad visas en varning när du exporterar till HTML om att befintliga BASIC-makron går förlorade.  
Utskriftslayout  
Markera här om även utskriftslayouten för det aktuella dokumentet ska exporteras.  
4.0 och MS Internet Explorer fr.o.m.  
Kopiera lokal grafik till Internet  
Om Du aktiverar detta alternativ så inkluderas inbäddad grafik med dokumentet vid uppladdning till vald Internet-server via FTP.  
Spara dokumentet via dialogrutan Spara som och ange en giltig fullständig URL på Internet som filnamn.  
HTML-filtret stödjer CSS2 (Cascading Style Sheets Level 2) för utskrift av dokument.  
Dessa funktioner är bara tillgängliga om export av utskriftslayout aktiveras.  
Teckenuppsättning  
Här väljer du en teckenuppsättning för exporten.  
Alternativ Textdokument  
Här kan du göra olika globala inställningar som definierar hur textdokument ska behandlas i %PRODUCTNAME.  
De här inställningarna gäller för alla nya %PRODUCTNAME Writer-dokument som du skapar.  
En del inställningar kan du även göra för det aktuella textdokumentet, om du sedan sparar det.  
De globala inställningarna sparas automatiskt.  
Standardteckensnitt (västliga)  
Med det här kommandot öppnar du en dialogruta där du ställer in standardteckensnitt.  
Standardteckensnitt (asiatiska)  
Om du har aktiverat stödet för asiatiska språk under Verktyg - Alternativ - Språkinställningar - Språk, ställer du in asiatiska standardteckensnitt här.  
Vy  
Här kan du göra förinställningar för visningen av vissa objekt i dokument och fönsterelement.  
Hjälplinjer  
I det här området visas visningsalternativ för begränsningar.  
Följande inställningar finns:  
Textbegränsningar  
Om den här rutan är aktiverad visas sidmarginalerna som tunna linjer.  
Tabellbegränsningar  
Om den här rutan är markerad inramas tabellceller av en tunn linje.  
Områdesbegränsningar  
Om den här rutan är markerad visas områdesbegränsningarna.  
Hjälplinjer vid förflyttning  
Det gör det lättare att placera ramen exakt i förhållande till linjalvärdena.  
Enkla handtag  
Om den här rutan är aktiverad så visas handtagen (de åtta punkterna i en begränsningsrektangel) som enkla kvadrater utan 3D-effekt.  
Stora handtag  
Om den här rutand är markerad så visas handtagen (de åtta punkterna i en begränsningsrektangel) större än vanligt.  
Vy  
Här kan du ställa in vilka rullningslister och linjaler som ska vara synliga.  
Horisontell rullningslist  
Här kan du dölja och visa den horisontella rullningslisten.  
Vertikal rullningslist  
Här kan du dölja och visa den vertikala rullningslisten.  
Horisontell linjal  
Här kan du dölja och visa den horisontella linjalen.  
Du väljer måttenhet i listrutan.  
Vertikal linjal  
Här visar och döljer du den vertikala linjalen.  
Du väljer måttenhet i listrutan.  
Mjuk rullning  
Här väljer du om sidan ska rullas mjukt.  
Hastigheten är beroende av vilken yta som ska rullas och vilket färgdjup som ska visas.  
Visa  
I det här området väljer du vilka dokumentelement som ska visas på bildskärmen.  
Grafik och objekt  
Om du markerar så visas grafik och objekt i dokumentet på bildskärmen.  
Om de är dolda så visas i stället tomma ramar som platshållare.  
Visningen av grafik kan du även styra via ikonen Grafik Grafik.  
Den här ikonen visas på verktygslisten om du har öppnat ett textdokument.  
När detta alternativ är avstängt laddas ingen grafik från Internet.  
När det finns grafiska objekt utan storleksangivelse i en tabell och någon besöker sidan, kan det uppstå problem med visningen av sidan om en äldre HTML-standard används.  
Tabeller  
Markera här om du vill att de tabeller som finns i dokumenten ska visas på bildskärmen.  
Teckningar och kontrollfält  
Markera här om teckningar och kontrollfält som finns i dokument ska visas på bildskärmen.  
Fältnamn  
Markera den här rutan om du vill att motsvarande fältkommando ska visas i ditt dokument i stället för innehållet i ett fält.  
När ett textdokument är öppet kan du även styra denna visning via menyn Visa - Fältkommandon Visa - Fältkommandon.  
Anteckningar  
Aktivera den här rutan om alla anteckningar och skript som finns i dina dokument ska visas som små rutor i färg.  
Om du vill läsa eller redigera innehållet dubbelklickar du på den önskade rutan.  
Bakgrund  
Vissa textelement kan med en grå bakgrund framhävas mot den vanliga texten.  
Dessa bakgrunder finns inte med på utskriften.  
I det här området kan Du definiera detta för följande element:  
Förteckningsposter (inte för HTML-dokument)  
Med detta alternativ förses infogade förteckningsposter förteckningsposter med en grå bakgrund.  
Förteckningar (inte för HTML-dokument)  
Om du markerar den här rutan visas infogade förteckningar förteckningar med grå bakgrund.  
Fotnoter (inte för HTML-dokument)  
Med detta alternativ förses fotnotsnummer fotnotsnummer med en grå bakgrund.  
Måttenhet (bara för HTML-dokument)  
Här väljer du måttenhet för HTML-dokument.  
Fält  
Med detta alternativ förses infogade fält fält med en grå bakgrund.  
Standardteckensnitt  
Med det här kommandot öppnas en dialogruta där du kan ställa in standardteckensnitt.  
Via de här inställningarna bestämmer du vilka standardteckensnitt som ska användas i de färdiga formatmallarna.  
Förutom standardteckensnitten kan du vid behov även ändra eller anpassa standardmallen för textformat.  
Standardteckensnitt  
Standard  
Här bestämmer Du vilket teckensnitt som ska användas i styckeformatmallen Standard.  
Eftersom nästan alla styckeformatmallar som medföljer programmet bygger hierarkiskt på styckeformatmallen Standard bestämmer Du härmed även teckensnittet för nästan alla färdiga styckeformatmallar i textområdet förutsatt att inte styckeformatmallen särskilt definierats med ett annat teckensnitt.  
Överskrift  
Här definierar Du standardteckensnittet i styckeformatmallarna för överskrifter och alla styckeformatmallar som baseras på dessa.  
För överskrifter lämpar sig främst sanserif-teckensnitt (utan seriffer) som t ex Arial Helvetica.  
Lista  
Det standardteckensnitt som definieras här används i styckeformatmallar för listor, numreringar och punktuppställningar och alla styckeformatmallar som baseras på dessa.  
De här styckeformatmallarna tilldelas automatiskt av programmet när ett numrerings - eller punktuppställningsstycke formateras via Format - Numrering / punktuppställning... Format - Numrering / punktuppställning...  
Bildtext  
Det standardteckensnitt som definieras här används i etiketter för bilder, tabeller och alla styckeformatmallar som baseras på dessa.  
Förteckning  
Det standardteckensnitt som definieras här används i styckeformatmallar för användardefinierade förteckningar, index, innehållsförteckningar och alla styckeformatmallar som baseras på dessa.  
Bara för det aktuella dokumentet  
Markera denna kryssruta om ändringarna i standardteckensnitten endast ska gälla för det aktuella dokumentet.  
Annars kommer ändringarna att gälla för alla nya dokument som skapas.  
Ändra standardmall  
Skriv ut  
Här kan du undanta vissa objekttyper från utskrift, välja utskrift av endast vänster - eller högersidor, definiera utskrift i omvänd ordningsföljd eller utskrift av prospekt.  
Dessutom väljer du var anteckningar ska skrivas ut, pappersmagasin och faxdrivrutin.  
De här inställningarna gäller sedan för alla textdokument som skrivs ut.  
Om du bara vill ändra inställningar för det aktuella dokumentet använder du kommandoknappen Fler i dialogrutan Arkiv - Skriv ut.  
Innehåll  
Här bestämmer du vilket dokumentinnehåll som ska skrivas ut.  
Du kan välja bland följande alternativ:  
Grafik  
Om den här rutan är markerad skrivs grafikobjekt i textdokument ut.  
Tabeller  
Om den här rutan är markerad skrivs tabeller i textdokument ut.  
Teckningar (inte för HTML-dokument)  
Om den här rutan är markerad skrivs grafik, som har skapats med ritfunktionerna, ut i textdokument.  
Kontrollfält  
Om rutan är markerad skrivs kontrollfält som infogats i textdokumentet ut.  
Bakgrund  
Om den här rutan är markerad skrivs bakgrunder som infogats i textdokument ut.  
Svart utskrift  
Markera den här rutan om text alltid ska skrivas ut i svart.  
Sidor  
I det här området anger du hur %PRODUCTNAME ska behandla flersidiga textdokument vid utskrift.  
Vänstersidor (inte för HTML-dokument)  
Om kryssrutan har markerats skrivs alla vänstersidor i dokumentet ut.  
Högersidor (inte för HTML-dokument)  
Om kryssrutan har markerats skrivs alla högersidor i dokumentet ut.  
Omvänt  
Om den här rutan är markerad skrivs dokument ut i omvänd ordningsföljd.  
Sista sidan i dokumentet skrivs då ut först.  
Då slipper du sortera sidorna efter utskrift.  
Prospekt  
Genom att markera den här kryssrutan kan du skriva ut dokumentet som prospekt.  
Då behandlar %PRODUCTNAME textdokument på följande sätt:  
Om du skriver ut ett dokument i stående format skrivs två motstående sidor i prospektet ut bredvid varandra.  
Om din skrivare klarar dubbelsidig utskrift kan du skapa ett färdigt prospekt utan att behöva sammanfoga sidorna efter utskrift.  
Om din skrivare bara klarar enkelsidig utskrift kan du uppnå samma effekt genom att först skriva ut alla förstasidor med alternativet Högersidor markerat och sedan lägga tillbaka hela pappersbunten i skrivaren igen och skriva ut på baksidorna med alternativet Vänstersidor markerat.  
Det enda du behöver se upp med är skrivarens utskriftsriktning.  
Anteckningar  
Inga  
När detta alternativ valts ignoreras anteckningar och skrivs inte ut.  
Endast anteckningar  
Om detta alternativ markeras skrivs alla anteckningar som gjorts för ett dokument ut.  
Själva dokumentet skrivs inte ut.  
Dokumentslut  
Om detta alternativ markerats skrivs dokumentsidorna ut först och sedan tillhörande anteckningar.  
Sidslut  
Om detta alternativ markerats skrivs dokumentet ut med anteckningarna nedtill på varje sida.  
Övrigt  
Skapa enstaka utskriftsjobb  
Om den här rutan är markerad börjar varje dokument som skrivs ut på ny sida även om du använder en skrivare med dubbelsidig utskrift.  
Annars kan t.ex. första sidan i andra satsen hamna på baksidan av det ark på vilket sista sidan i första satsen skrivits ut.  
Pappersmagasin från skrivarinställning  
Via detta alternativ anger du, för skrivare med flera pappersmagasin, om pappersmagasin ska väljas från skrivarens systeminställningar.  
Fax  
Om du har ett faxprogram installerat på din dator och vill faxa direkt från textdokument ska du välja faxen i det här kombinationsfältet.  
Tabell  
Här definierar du egenskaper för tabeller i textdokument.  
Här gör du förinställningar för det inbördes förhållandet mellan kolumner och rader och för valt tabelläge.  
Dessutom kan du definiera de standardvärden som används när du flyttar / infogar kolumner och rader.  
Det finns mer information om detta i %PRODUCTNAME Writer - hjälpen under Anpassa tabell rubriken "Anpassa tabell".  
Standard  
Här gör du förinställningar för alla nya texttabeller som skapas i textdokument.  
Överskrift  
Markera den här rutan om den första raden i tabellen ska formateras med styckeformatmallen "Tabellöverskrift".  
Upprepa på varje sida  
Om en tabell måste delas upp på flera sidor och du vill att tabellöverskriften ska upprepas på varje sida markerar du den här rutan.  
Dela inte (inte för HTML)  
Om den här kryssrutan är markerad, kan tabellen inte delas vid sidbrytning.  
Du kan även göra den här inställningen via menykommandot Format - Tabell - Textflöde.  
Inramning  
Här kan du ställa in om tabellcellerna ska ha ramar som standard.  
Inmatning i tabeller  
Taligenkänning  
Om den här rutan är markerad känns tal igen som tal i en texttabell.  
Talen formateras i talformat.  
Du kan påverka hur justeringen görs med rutan Justering.  
Om rutan Taligenkänning inte är markerad, sparas tal i textformat och vänsterjusteras automatiskt liksom den text som skrivs in.  
Talformatsigenkänning  
Om den här rutan inte är markerad, godtas en inmatning bara om den görs i det format som har angetts för cellen i fråga.  
Andra inmatningar återställer formatet till Text.  
Om talformatet för cellen är inställt på t.ex. "-123,45 €", identifieras även inmatningar i formaten 123 eller 123 €som tal.  
Men om du skriver 1.1, tolkas detta som ett datum, vilket inte stämmer med det format som har angetts för cellen.  
Inmatningen formateras därför som text.  
Justering  
Om den här rutan är markerad högerjusteras tal alltid nere i cellen.  
Om den här rutan inte är markerad vänsterjusteras alltid tal uppe i cellen.  
Direkta formateringar påverkas inte av rutan Justering.  
Om du centrerar cellinnehåll direkt, förblir det centrerat, oavsett om det rör sig om text eller om tal.  
Flytta  
Här definierar du standardinställningar som gäller när rader och kolumner flyttas med hjälp av tangentbordet.  
Tryck samtidigt på Alt och en piltangent.  
Rad  
I det här rotationsfältet anger du ett värde för hur mycket raden ska flyttas.  
Kolumn  
I det här rotationsfältet anger du ett värde för hur mycket kolumnen ska flyttas.  
Infoga  
Här definierar du standardinställningar som gäller när fler rader och kolumner infogas med hjälp av tangentbordet.  
Tryck på Alt+Insert och sedan på en piltangent.  
Rad  
I det här rotationsfältet anger Du ett värde som ska användas som standardvärde för infogning av rader.  
Kolumn  
I det här rotationsfältet anger Du ett värde som ska användas som standardvärde för infogning av kolumner.  
Effekt av ändringar  
Här väljer Du hur spalter och rader ska påverka varandra och omgivningen eller hur hela tabellen ska påverkas.  
Fast  
Klicka här om Du vill att ändringar i en rad och / eller kolumn endast ska påverka den närmaste omgivningen.  
Den här inställningen kan Du även göra via ikonen Tabell: fast Tabell: fast, som visas i objektlisten när ett textdokument är öppet och markören står i en tabell.  
Fast, proportionell  
Klicka här om Du vill att ändringar i en kolumn och / eller rad ska påverka hela tabellen.  
På motsvarande sätt använder Du ikonen Tabell: fast, proportionell Tabell: fast, proportionell, som visas i objektlisten när ett textdokument är öppet och en tabell är markerad.  
Variabel  
Klicka här om Du vill att ändringar i en rad och / eller kolumn ska påverka tabellstorleken.  
När ett textdokument är öppet kan de olika lägena även ställas in via motsvarande ikon ikon i tabellobjektlisten.  
Formateringshjälp  
Här gör du inställningar för visningen av vissa tecken och för direktmarkören.  
En del av de här inställningarna kan du även göra för HTML-dokument.  
Visa  
I det här området definierar du vilka av de icke utskrivbara tecknen som ska visas på bildskärmen.  
Om du klickar på ikonen Kontrolltecken på / av Kontrolltecken på / av på verktygslisten visas alla tecken som du har markerat här i dokumentet.  
Stycketecken  
Om du markerar den här rutan visas stycketecken.  
Stycketecknet innehåller även formatinformation för ett stycke.  
Användardefinierade bindestreck  
Om du markerar den här rutan visas användardefinierade bindestreck.  
Detta är dolda bindestreck som du kan mata in inuti ett ord med Kommando+" - "Ctrl+" -".  
I slutet av raden avstavas det här ordet bara på ett ställe där ett användardefinierat bindestreck har matats in oavsett om den automatiska avstavningen är aktiverad eller inte.  
Blanksteg  
Om du markerar den här rutan, så markeras varje blanksteg i texten med en liten punkt.  
Fast mellanrum  
Om du markerar den här rutan visas fasta mellanrum som gråa rutor.  
Du infogar fast mellanrum med tangentkombinationen Kommando+Blanksteg Ctrl+Blanksteg.  
Tabulatorer  
Markera den här rutan om du vill att tabbarna ska visas som tecken.  
Brytningar  
Om den här kryssrutan är markerad så visas de radslut som har infogats med Skift+Retur.  
Dessa brytningar anger ett tvingande radbyte utan att ett nytt stycke påbörjas.  
Dold text (inte för HTML-dokument)  
När du har infogat text med fältfunktionerna Villkorlig text eller Dold text kan du med den här kryssrutan bestämma om den här texten ska visas eller döljas.  
Dolda stycken (inte för HTML-dokument)  
När du har infogat text med fältfunktionen Dolt stycke kan du med den här kryssrutan bestämma om texten ska visas eller döljas.  
Den här kryssrutan har samma funktion som menykommandot Visa - Dolda stycken Visa - Dolda stycken som är tillgängligt när ett textdokument är öppet.  
Direktmarkör (inte för HTML-dokument)  
I det här området ställs direktmarkörens samtliga egenskaper in.  
Direktmarkör  
Om Du markerar den här kryssrutan aktiveras direktmarkören.  
Du har tillgång till samma funktion via ikonen Direktmarkör Direktmarkör på verktygslisten, när ett textdokument är öppet.  
Infoga (inte för HTML-dokument)  
Här definierar Du direktmarkörens infogningsalternativ.  
Om du klickar med direktmarkören på en plats i dokumentet, infogas där ett stycke som, beroende på vilket alternativ Du har valt, kan ha olika egenskaper.  
Du kan välja mellan följande alternativ:  
Styckejustering  
När du använder direktmarkören justeras stycket.  
Beroende på var du klickar med musen vänsterjusteras, centreras eller högerjusteras stycket.  
Innan du klickar visar markören med en triangel vilken justering som är inställd.  
Vänster styckemarginal  
När du använder direktmarkören sätts det vänstra styckeindraget vid den horisontella position där du klickar med direktmarkören.  
Stycket vänsterjusteras.  
Tabulator  
När du använder direktmarkören infogas så många tabbar i det nya stycket som det behövs för att komma till den position där du klickar.  
Tabulator och blanksteg  
När du använder direktmarkören infogas så många tabbar och blanksteg i det nya stycket som det behövs för att komma till den position där du klickar.  
Samtliga infogningsalternativ gäller bara det aktuella stycke som skapas med direktmarkören.  
Färg  
I det här kombinationsfältet väljer Du färg för direktmarkören.  
Tillåt markör i skyddade områden  
Om du markerar den här rutan, kan Du placera markören i ett skyddat område men inte göra några ändringar.  
Ändringar  
Här definierar du om registrerade ändringar i dokumentet ska framhävas.  
Om du vill registrera eller visa ändringar väljer du menykommandot Redigera - Ändringar nÃ¤r du har Ã¶ppnat ett text - eller tabelldokument.  
Textvisning  
Här ställer du in visningen av de registrerade ändringarna.  
Med alternativfälten bestämmer du för vilken typ av ändringar vilket attribut och vilken färg ska användas för visning.  
I ett förhandsvisningsfält ser du hur den valda visningen ser ut.  
Infoga / Attribut  
Med detta alternativ definierar Du hur ny text som infogas i dokumentet ska visas.  
Radera / Attribut  
Med det här alternativet bestämmer du hur ändringar ska visas i dokumentet när en text har raderats.  
När du registrerar radering av en text, raderas texten inte utan förses med det valda attributet, t.ex. en genomstrykning.  
Attributändring / Attribut  
Med detta alternativ definierar Du hur ändringar av teckenattribut i ett dokument ska visas.  
Sådana ändringar omfattar t ex tilldelning av attributen Fet, Kursiv och Understrykning.  
Färg  
Här väljer du vilken färg som ska visas för ändringen.  
Färgen varierar beroende på vilken författare som har gjort ändringarna.  
Ändrade rader  
Markeringen kan infogas antingen i vänster - eller högermarginalen.  
Markering  
Här definierar du om och var ändrade rader i dokumentet ska markeras.  
Du kan också låta placeringen vara beroende av om det är en höger - eller en vänstersida och i så fall att markeringen alltid ska göras i den utvändiga eller invändiga marginalen.  
Färg  
Här väljer Du färg på markeringen för ändrade rader.  
Bildtext  
I den här dialogrutan kan du göra bildtextinställningar för valda objekttyper.  
Bildtext  
Klicka på rutan framför den objekttyp som bildtextinställningarna ska gälla för.  
Inställningar  
I det här området gör du de inställningar som bara ska gälla för den valda objekttypen.  
Alternativen motsvarar dem på menyn Infoga - Bildtext....  
Nedanför listrutorna visas objektets beteckning inklusive numreringstyp.  
Kategori  
Här visas det markerade objektets kategori.  
Objektnamnet kan du ändra vid behov.  
Du kan också välja en annan kategori i listrutan.  
I %PRODUCTNAME används Illustration, Tabell och Text som standardkategorier.  
Numrering  
Här väljer du vilken typ av numrering som du vill ha.  
Bildtext  
I den här listrutan skriver du bildtexten.  
Position  
I den här listrutan anger du om bildtexten ska placeras ovanför eller nedanför objektet.  
Nivå  
Här väljer du den överskrifts - respektive kapitelnivå vid vilken numreringen ska börja om när nivån ändras.  
Skiljetecken  
Ange här det tecken som direkt ska följa efter numret på rubrik - respektive kapitelnivå.  
Allmänt  
Här gör du allmänna inställningar för textdokument.  
Uppdatera länkar vid laddning  
Alltid  
Med det här alternativet uppdateras länkar automatiskt när ett dokument laddas.  
På begäran  
Med detta alternativ uppdateras länkar bara på begäran när ett dokument laddas.  
Aldrig  
Med detta alternativ uppdateras länkar inte automatiskt när ett dokument laddas.  
Fält och diagram  
Fältkommandon automatiskt  
Markera den här rutan om fältkommandon som finns i dokumenten ska uppdateras automatiskt.  
Uppdatera diagram automatiskt  
Diagram uppdateras automatiskt om du markerar den här rutan.  
Kryssrutan går bara att använda om Fältkommandon automatiskt är markerad.  
Bildtext  
Här anger Du hur de beskrivningar ska se ut som ges till de tabeller, bilder och ramar som infogas i textdokument och de %PRODUCTNAME -objekt som infogas som OLE-objekt.  
Automatiskt  
Om du markerar den här rutan formateras objekten som har valts i Objekturval automatiskt enligt reglerna som har definierats där.  
Om inga regler för objekt är definierade där rättar sig bildtexten till ett infogat objekt efter de definierade inställningarna på menyn Infoga - Bildtext  
Objekturval  
...  
Med den här kommandoknappen öppnar du dialogrutan Bildtext där du kan göra förinställningar för enskilda dokumenttyper.  
Måttenhet  
Här väljer du måttenhet för textdokument.  
Tabulatoravstånd  
I detta rotationsfält anger Du vilket avstånd de enskilda tabbarna ska ha.  
Det avstånd som Du väljer visas på den horisontella linjalen.  
Kompatibilitet  
I de olika ordbehandlingsprogrammen är formateringsdefinitionerna inte identiska.  
När Du skapar dokument med %PRODUCTNAME Writer och de ändå ska vara kompatibla framför allt till MS Word, så kan Du ställa in detta här.  
Inställningarna i detta område kan bara göras för ett aktuellt dokument och gäller också bara för detta.  
Kryssrutorna är därför bara tillgängliga om det finns ett öppnat textdokument.  
Addera alla stycke - och tabellavstånd i det aktuella dokumentet  
I %PRODUCTNAME Writer är styckeavstånd definierade på annat sätt än i MS Word-dokument.  
Om du har ställt in ett övre och ett nedre avstånd mellan två stycken, så adderas dessa för MS Word-dokument, medan %PRODUCTNAME Writer tar det större av de båda.  
Markera den här rutan om avstånden mellan stycken och mellan tabeller ska adderas i %PRODUCTNAME Writer.  
Lägg till stycke - och tabellavstånd vid början av sidor  
Om denna ruta är markerad så beaktas styckeavståndet uppåt också i början på en sida eller kolumn även när stycket finns på dokumentets första sida.  
Samma sak gäller vid en sidbrytning.  
När Du importerar ett MS Word-dokument så adderas avstånden automatiskt vid konverteringen.  
Justera tabulatorposition  
Om den här rutan är markerad formateras centrerade och högerjusterade stycken som innehåller tabbar helt och hållet centrerat eller högerjusterat.  
Om rutan är markerad, högerjusteras t.ex. bara texten till höger om den sista tabulatorn, medan texten till vänster stannar kvar på sin plats.  
Alternativ - HTML-dokument  
Här gör du grundinställningar för %PRODUCTNAME -dokument i HTML-format.  
Du väljer bl.a. vad som ska visas på bildskärmen eller på utskriften, om sidorna på bildskärmen ska rullas mjukt eller i vilka färger nyckelorden i källtexterna ska visas.  
Raster  
Här ställer du in att att sidorna i dokument ska ha ett justerbart raster.  
Om du vill kan du synkronisera det "magnetiska" stödrastret med det här rastret.  
Raster  
I det här området bestämmer du vilken indelning rastret ska ha.  
Du kan använda olika måttenheter.  
Använd stödraster  
Om du klickar här kan ramar, teckningselement och formulärfunktioner bara flyttas mellan olika rasterpunkter.  
Om du flyttar ett objekt och håller ner Kommandotangenten Ctrl-tangenten ändras stödrastrets status medan du flyttar.  
Synligt raster  
Med det här kommandot visas rastret.  
Den här funktionen finns även som ikon på alternativlisten i ett öppet presentationsdokument. ikon på alternativlisten i ett öppet teckningsdokument. ikon med namnet Visa raster på alternativlisten om ett formulärobjekt är markerat.  
Du kan även ange om rastret ska var synligt eller inte med alternativet Raster synligt på sidans snabbmeny.  
Dessutom kan Du med kommandot Raster främst på snabbmenyn ange om rastret ska ligga framför eller bakom objekt.  
Du kan även ange om rastret ska var synligt eller inte med kommandot Raster synligt på sidans snabbmeny.  
Dessutom kan du med kommandot Raster främst på snabbmenyn ange om rastret ska ligga framför eller bakom objekt.  
Horisontell upplösning  
Här definierar du avståndet mellan rasterpunkter på X-axeln i önskad måttenhet.  
Horisontell indelning  
Här anger Du antalet mellansteg mellan rasterpunkterna på X-axeln.  
Därigenom kan Du finfördela rasterindelningen ytterligare.  
Vertikal upplösning  
Här anger Du avståndet mellan rasterpunkterna på Y-axeln i önskad måttenhet.  
Vertikal indelning  
Här anger Du antalet steg mellan rasterpunkterna på Y-axeln.  
Därigenom kan Du finfördela rasterindelningen ytterligare.  
Synkronisera axlar  
Markera den här kryssrutan om Du vill ändra de aktuella rasterinställningarna symmetriskt.  
Upplösningen och indelningen för X - och Y-axeln är då alltid lika.  
På sidans snabbmeny finns ytterligare kommandon:  
På sidans snabbmeny finns ytterligare kommandon:  
Raster främst Raster främst  
Med det här alternativet placerar Du det synliga rastret framför alla objekt.  
Med det här alternativet placerar Du det synliga rastret framför alla objekt.  
Hjälplinjer främst Hjälplinjer främst  
Med det här alternativet visar Du hjälplinjerna framför alla objekt.  
Med det här alternativet visar Du hjälplinjerna framför alla objekt.  
Källtext  
Här bestämmer du med vilken färg kända och okända textsegment ska visas i källtextredigeraren.  
Färgtilldelning för syntaxframhävning  
Välj färg för de olika textelementen i listrutorna.  
SGML  
Här väljer du färg för de taggar i det sidbeskrivande språket SGML som inte hör till HTML-standard.  
I normala HTML-dokument är det den första raden.  
Kommentar  
Här väljer du färg för kommentarer i källtexten.  
Nyckelord  
Här väljer du färg för nyckelord.  
Okänd  
Här väljer du färg för alla övriga textelement.  
Bakgrund  
I den här dialogrutan väljer du bakgrund för HTML-dokument.  
Bakgrund gäller för nya HTML-dokument och för sådana som du laddar om de inte har definierat en egen bakgrund.  
Mer information  
Alternativ Tabelldokument  
Du bestämmer bland annat vilket innehåll som ska synas och i vilken riktning markören flyttas när du har matat in data i en cell.  
Du definierar sorteringslistor, bestämmer det generella antalet decimaler för visningen och förinställningar för hur ändringar registreras och framhävs.  
En del inställningar gäller bara globalt om det aktiva dokumentet inte är ett dokument av den här typen.  
Om ett dokument av den här typen är aktivt, gäller en del inställningar bara för det aktuella dokumentet och sparas med det.  
Vy  
Här bestämmer du vilka element i huvudfönstret som ska visas och om värdena i tabellen ska framhävas.  
Optisk hjälp  
Här definierar du vilka linjer som ska visas.  
Gitterlinjer  
Markera här om du vill att gitterlinjerna mellan cellerna ska visas på bildskärmen.  
När det gäller utskrift gör du motsvarande inställning under Format - Sida - fliken Tabell med rutan Tabellgitter.  
Färg  
I den här listrutan väljer du färg för de visade gitterlinjerna.  
Sidbrytningar  
Om du aktiverar den här kryssrutan, visas sidbrytningarna för ett definierat utskriftsområde.  
Hjälplinjer när objekt flyttas  
Markera den här rutan om hjälplinjer ska visas när du flyttar teckningar, ramar, grafikobjekt och andra objekt.  
De här linjerna hjälper dig att justera objekt.  
Enkla handtag  
Om den här rutan är markerad, visas handtagen (de åtta punkterna i en begränsningsrektangel) som enkla kvadrater utan 3D-effekt.  
Stora handtag  
Om den här rutan är markerad, visas handtagen (de åtta punkterna i en begränsningsrektangel) större än normalt.  
Visa  
I det här området väljer du vad som ska visas på bildskärmen.  
Formler  
Markera den här rutan om du vill att formlerna ska visas i cellerna i stället för resultaten.  
Nollvärden  
Markera här om du vill att tal med värdet 0 ska visas.  
Anteckningsmarkör  
Markera här om du vill att anteckningar i cellerna ska visas.  
En liten rektangel i det övre högra hörnet i en cell visar att det finns en anteckning.  
De här rektanglarna aktiverar du under Verktyg - Alternativ - Tabelldokument - Vy genom att markera rutan Anteckningsmarkör.  
På snabbmenyn till en cell som innehåller en anteckning hittar du kommandot Visa anteckning.  
När du klickar på det här kommandot visas anteckningen till den här cellen hela tiden och kommandot bockmarkeras.  
Du infogar och redigerar anteckningar med menykommandot Infoga - Anteckning.  
De anteckningar som alltid visas kan Du klicka på och redigera direkt.  
Genom att dubbelklicka på en anteckning flyttar Du cellmarkören till motsvarande cell.  
Framhäv värden  
Markera denna ruta om alla värden i tabellen ska framhävas i färg.  
Textceller formateras med svart färg, celler som innehåller tal är blå och andra celler (formler, logiska värden, datum etc.) är gröna.  
När detta kommando är aktivt visas inte de färger som har angetts i dokumentet.  
Färgerna finns dock kvar och visas igen när Du avmarkerar kryssrutan.  
Ankare  
När du markerar den här rutan visas ankarsymbolen för ett markerat grafiskt objekt i ett dokument.  
Textspill  
Den indikerar att texten fortsätter.  
Om den här rutan inte är markerad visas inte triangeln.  
Visa referenser i färg  
Om Du tar bort markeringen visas referenserna i formlerna från inmatningsraden inte längre i färg.  
Om Du har markerat rutan ser Du varje enskild referens, t ex i form av "=B1:C2+D5:G9" både framhävd i färg i formler och i samma färg som cellområdets inramning, så snart Du markerar en cell som innehåller referensen för redigering.  
Objekt  
I detta område kan Du för tre objektgrupper definiera om de ska visas, döljas eller ersättas av platshållare.  
Objekt / grafik  
Här väljer Du om objekt och grafik ska visas, döljas eller ersättas av platshållare.  
Diagram  
Här väljer Du om diagram ska visas, döljas eller ersättas av platshållare.  
Ritobjekt  
Här väljer Du om ritobjekt ska visas, döljas eller ersättas av platshållare.  
Fönster  
I det här området anger Du för några hjälpelement om de ska visas i tabellen eller ej.  
Kolumn - och radhuvuden  
Markera den här rutan om Du vill att kolumn - och radhuvuden ska visas.  
Horisontell rullningslist  
Markera den här rutan om Du vill att en rullningslist för horisontell förflyttning av stora tabeller ska visas vid tabellfönstrets nedre ram.  
Vertikal rullningslist  
Markera den här rutan om Du vill att en rullningslist för vertikal förflyttning av stora tabeller ska visas vid tabellfönstrets högra ram.  
Tabellflik  
Markera den här rutan om Du vill att tabellflikar ska visas vid tabellernas nedre ram så att man kan växla mellan visade tabeller.  
Om Du har inaktiverat den här hjälpen, kan Du bara skifta mellan tabellerna via Navigator.  
Om Du aktiverar tabellregistren igen efter inaktiveringen, gäller det bara för de nya dokument som skapats eller laddats.  
Dispositionssymboler  
Här markerar Du om Du vill se dispositionsssymbolerna i kanten av tabellen, såvida Du har definierat en disposition.  
Allmänt  
Här bestämmer bl.a. du vad som händer när du trycker på returtangenten i en tabell.  
Metriker  
Måttenhet  
Här väljer du måttenhet i tabeller.  
Tabulatoravstånd  
Ange tabulatoravståndet i det här rotationsfältet.  
Inmatningsinställningar  
Tryck Retur för att flytta markering  
Om du klickar på det här fältet och t.ex. väljer till höger i listrutan bredvid, markeras nästa cell till höger när du trycker på returtangenten.  
Retur växlar till redigeringsläge  
Med denna funktion kan Du redigera den markerade cellen direkt efter att Du tryckt på returtangenten.  
Utöka formatering  
Med den här funktionen överförs formateringarna för en cell automatiskt till de angränsande tomma cellerna.  
Om du t.ex. har formaterat cellinnehållet med fetstil, kommer alla värden som du matar in i tomma celler i samma område också att ha fetstil.  
Celler som redan är formaterade ändras inte.  
Om du använder tangentkombinationen Kommando Ctrl +* [multiplikationstecknet på den numeriska delen av tangentbordet] ser du området som påverkas av den här funktionen.  
Alla värden som du matar in i det här området får den definierade formateringen.  
När du sätter markören i en cell utanför området gäller standardformateringen igen.  
Utöka referenser i kanterna när kolumner / rader infogas  
Slå på denna funktion om referenser vid infogning av rader eller kolumner ska utökas direkt bredvid / över / under referensområdet.  
Detta sker endast om den tidigare referensen har en utbredning som omfattar minst två celler i den riktning som infogningen har gjorts.  
Exempel:  
Om Du refererar till en formel i området A1:B1 och Du infogar en ny kolumn efter kolumn B, så utökas referensen till A1:C1 om Du har markerat denna ruta.  
Om Du refererar till området A1:B1 och infogar en ny rad under rad 1, utökas referensen inte eftersom det bara finns en enda cell i den lodräta riktningen.  
Om Du infogar rader eller kolumner i mitten av ett referensområde utökas referensen självklart alltid.  
Framhäv markering i kolumn - / radhuvuden  
Om den här rutan är markerad framhävs markerade kolumner och rader i kolumn - och radhuvudena.  
Använd skrivarmått för textformatering  
Om den här rutan är markerad används skrivarmåtten inte bara för utskrift utan även för formatering av visningen på bildskärmen.  
Sorteringslistor  
Här visas alla användardefinierade listor.  
Vidare kan du själv definiera och redigera listor.  
Listor  
Här visas alla tillgängliga listor och du kan välja en för redigering.  
Poster  
Här ser du innehållet i den markerade listan och kan redigera det.  
Kopiera lista från  
I det här fältet kan Du definiera från vilken tabell och vilka celler en lista ska kopieras och tilldela den området Listor.  
Det i tabellen markerade området är här förinställt.  
Kopiera  
Med den här kommandoknappen kopierar Du innehållet i de celler som anges i Kopiera lista från.  
Om Du har markerat en referens av sammanhängande rader och kolumner efter att ha klickat på kommandoknappen, visas dialogrutan Kopiera lista där Du kan ange om referensen ska sorteras radvis eller kolumnvis till sorteringslistor.  
Nytt / Ignorera  
Om du vill skapa en ny lista, kan du klicka på den här kommandoknappen och mata in den här listans innehåll i området Poster.  
Kommandoknappen ändrar sin funktion från Nytt till Ignorera.  
Du kan ta bort den lista du nyss skapat med kommandoknappen Ignorera.  
Lägg till / Ändra  
Med den här kommandoknappen kan Du överta den nya listan i området Listor.  
Om Du i området Poster skulle göra ändringar i redan befintliga listor, skiftar kommandoknappen funktion från Lägg till till Ändra och Du kan överta den ändrade listan genom att klicka på Ändra.  
Kopiera lista  
Här kan du kopiera de markerade cellerna till en sorteringslista.  
Lista från  
Vid kopiering ignoreras celler utan text.  
Rader  
Markera detta alternativfält om Du vill sammanfatta innehållet i de markerade raderna i en lista.  
Kolumner  
Markera detta alternativfält om Du vill sammanfatta innehållet i de markerade kolumnerna i en lista.  
Beräkna  
Här kan du göra förinställningar för tabellberäkningar.  
Du definierar hur %PRODUCTNAME Calc ska reagera vid cirkulära referenser i tabelldokument, ställer in basen för datumangivelser och antalet decimaler samt anger om programmet ska ta hänsyn till versaler / gemener vid tabelljämförelser.  
Cirkulära referenser  
I det här området kan du begränsa det antal approximeringssteg som ska utföras vid iterativa beräkningar.  
Vidare kan du fastställa med vilken noggrannhet som resultaten ska anges.  
Iterationer  
Markera den här rutan om %PRODUCTNAME Calc ska försöka beräkna ett resultat för tabelldokument med cirkulära referenser (referenser till sig själv) med hjälp av upprepade beräkningssteg.  
Om den här rutan inte är markerad, vilket är förinställningen, leder en cirkulär referens i tabellen till ett felmeddelande (vilket är rimligt, eftersom cirkulära referenser oftast inte är önskvärda utan uppstår genom misstag).  
Exempel:  
Du vill dela upp ett försäljningspris i nettopris och mervärdesskatt (moms).  
Därför skriver du t.ex. i A5 texten "FP", i A6 texten "Netto" och i A7 texten "Moms ".  
Mata nu in försäljningspriset (t.ex. 100) i B5.  
I cell B6 ska nettopriset stå och i B7 mervärdesskatten.  
Du vet att momsen räknas ut som "nettopriset gånger 25%" och att nettopriset returneras när du drar momsen från försäljningspriset.  
Alltså skriver du i B6 formeln "=B5-B7" för nettopriset, och i cell B7 skriver du formeln "=B6*0,25 "för momsen.  
Om iterationen är avstängd, får du följande felmeddelande på statuslisten: "Cirkulär referens".  
Om du aktiverar iterationen beräknas formlerna korrekt.  
A  
B  
5  
FP  
100  
6  
Netto  
=B5-B7  
7  
Moms  
=B6*0,25  
Steg  
Här anger du det största tillåtna antalet iterationssteg i beräkningen.  
Minsta ändringsvärde  
Om skillnaden underskrider detta värde avbryts iterationen.  
Datum  
I det här området väljer du startdatum för den interna omvandlingen av dagar till tal.  
1899-12-30 (standard)  
Som standard tilldelas datumet 1899-12-30 numret noll.  
1900-01-01 (StarCalc 1.0)  
Här väljer du att datumet 1 januari 1900 ska vara dag nummer noll.  
Välj den här inställningen om du öppnar en tabell som är skapad i StarCalc 1.0 och innehåller datumangivelser.  
1904-01-01  
Här väljer du att datumet 1 januari 1904 ska vara dag nummer noll.  
Den här inställningen gäller för vissa importformat i externa tabeller.  
Versalkänslig  
Om du markerar den här rutan, kommer stora och små bokstäver att betraktas som olika tecken vid jämförelse av cellinnehåll.  
Exempel:  
Skriv texten "Test" i cell A1 och texten "test "i cell B1.  
Skriv sedan formeln "=A1=B1" i cell C1.  
I annat fall skulle resultatet bli SANT.  
Textfunktionen IDENTISK tar alltid hänsyn till skillnaden mellan stor och liten bokstav oavsett vilken inställning du gör i den här dialogrutan.  
Antal decimaler  
Här bestämmer du hur många decimaler som ska visas i decimaltal som har formaterats med formatet Standard.  
Talen visas avrundade men sparas utan avrundning.  
Precision som visat  
Om du markerar den här rutan, fortsätter beräkningen med värden avrundade enligt den regel som du har angett.  
Diagram representeras med angivna värden.  
Om rutan inte är markerad, avrundas visningen till t.ex. två decimaler medan beräkningarna internt görs med alla decimaler.  
Sökkriterier = och < > måste matcha hela celler  
Om den här kryssrutan är markerad, måste de sökkriterier som du har valt för databasfunktionerna exakt stämma med hela cellen.  
Om den här rutan är markerad, beter sig %PRODUCTNAME Calc precis som MS Excel vid sökningar i celler i databasfunktionerna.  
.* på följande plats:  
Inverkan på sökningen:  
win  
"win" hittas; däremot inte "win95 "eller "windows"  
win.*  
"win" och "win95 "hittas; däremot inte "OS2win"  
.*win  
"win" och "OS2win "hittas; däremot inte "win95" eller "windows "  
.*win.*  
"win", "win95", "OS2win" och "windows "hittas  
Om den här kryssrutan inte är markerad, fungerar sökordet "win" på samma sätt som ".*win* ", d.v.s. det räcker om sökordet finns någonstans inuti cellen vid en sökning i databasfunktionerna.  
Tillåt reguljära uttryck i formler  
Om den här rutan är markerad går det att använda reguljära uttryck vid sökning och jämförelse av strängar.  
Detta gäller t.ex. databasfunktionerna, LETARAD, LETAKOLUMN och SÖK.  
Sök kolumn - / radetiketter automatiskt  
Om du markerar den här kryssrutan kan du använda texten i en cell till att peka på kolumnområdet nedanför texten eller på radområdet till höger om texten.  
Texten måste bestå av minst ett ord och får inte innehålla någon operator.  
Exempel: i cell E5 står texten "Europa".  
Under den i cell E6 står värdet 100 och i cell E7 värdet 200.  
Om den här rutan är markerad kan du nu skriva formeln: =SUMMA( Europa) i cell A1.  
Ändringar  
Här finns alternativ som du kan använda om du vill att registrerade ändringar i ditt dokument ska visas i färg.  
Om du vill registrera ändringar i arbetet, väljer du Redigera - Ändringar.  
Färggivning för ändringar  
I detta område definierar Du de önskade färgerna för fyra olika ändringar i dokumentet.  
Med posten "Efter författare" bestäms färgen automatiskt av %PRODUCTNAME och varieras med hänsyn till den författare som gör ändringarna.  
Ändringar  
Här kan Du bestämma en färg för ändringar av cellinnehåll.  
Raderingar  
Ifall raderingar ska markeras med färger, väljer Du i detta kombinationsfält en färg.  
Infogningar  
Ifall infogningar ska markeras med färger, väljer Du i detta fält en färg.  
Förskjutningar  
Ifall förskjutning av innehåll ska markeras med färger, väljer Du i detta fält en färg.  
Skriv ut  
Här gör du utskriftsinställningar för tabelldokument.  
Om du vill göra inställningar för det aktuella dokumentet väljer du Arkiv - Skriv ut, kommandoknapp Fler.  
Om du vill göra förinställningar för alla tabelldokument väljer du Verktyg - Alternativ - Tabelldokument - Skriv ut.  
Sidor  
Undertryck utmatning av tomma sidor  
Om den här rutan är markerad skrivs tomma sidor, som inte innehåller något cellinnehåll och inte något ritobjekt, inte ut.  
Cellattribut som kanter eller bakgrundsfärg är inget cellinnehåll.  
De tomma sidorna räknas inte med vid sidnumrering.  
Tabeller  
Skriv bara ut markerade tabeller  
Om den här rutan är markerad skrivs bara de markerade tabellerna ut, även om du väljer utskriftsområdet "Allt" i dialogrutan Arkiv - Skriv ut.  
Om du har matat in flera "sidor" som utskriftsområdet i dialogrutan Arkiv - Skriv ut skrivs bara de sidor (tabeller) ut som är markerade i utskriftsområdet.  
Om du vill markera en tabell håller du ner Ctrl-tangenten och klickar på tabellnamnet i undre kanten av arbetsområdet.  
Alternativ Presentation  
Här gör du inställningar för alla nya presentationsdokument.  
Bland annat bestämmer du vilket innehåll som ska visas på sidorna, vilken måttenhet som gäller, om och hur en justering mot rastret ska ske och om du vill att anteckningar och flygblad ska skrivas ut.  
Vy  
Här kan du välja mellan olika ersättningsvisningar.  
Genom att välja en ersättningsvisning påskyndar du uppdateringen av bildskärmen vid redigering.  
Ersättningsvisning  
För mycket komplicerade teckningselement tar det lite längre tid att uppdatera bildskärmen.  
Däremot visas den inte på bildskärmen.  
Antyd extern grafik  
Välj det här alternativet om bara konturerna av infogade grafikobjekt ska visas.  
När ett presentations - eller teckningsdokument är öppet kan du också nå den här funktionen med hjälp av ikonen ikonen ikonen med samma namn på alternativlisten.  
Konturläge  
Med den här rutan bestämmer du att bara konturen visas av fyllda teckningselement.  
Ytfyllningen visas inte.  
När ett presentations - eller teckningsdokument är öppet kan Du också ställa in konturläget med hjälp av ikonen Konturläge Konturläge Konturläge på alternativlisten.  
Antyd text  
Markera den här rutan om du vill att textfönster ska visas utan textinnehåll.  
Uppdateringen av bildskärmen går betydligt snabbare.  
När ett presentations - eller teckningsdokument är öppet kan du också nå den här funktionen med hjälp av ikonen ikonen ikonen med samma namn på alternativlisten.  
Visa bara fina linjer  
Om du markerar den här rutan visas linjer och inramningar bara som tunna linjer.  
Visningen är oberoende av den verkliga linjebredden.  
När ett presentations - eller teckningsdokument är öppet kan du också nå den här funktionen med hjälp av ikonen ikonen ikonen med samma namn på alternativlisten.  
Visa  
Linjaler synliga  
Markera den här rutan om du vill få tillgång till hjälplinjalerna med måttangivelser till vänster och ovanför arbetsområdet.  
Hjälplinjer vid förflyttning  
Markera den här rutan om du vill att hjälplinjer ska visas när du flyttar ett objekt.  
I %PRODUCTNAME skapas streckade hjälplinjer som förlänger sidorna på begränsningsrektangeln runt det markerade objektet så att den omfattar hela arbetsområdet.  
Detta gör det enklare att placera objekt.  
När ett presentations - eller teckningsdokument är öppet kan du också ställa in den här funktionen med hjälp av ikonen ikonen ikonen med samma namn på alternativlisten.  
Alla kontrollpunkter i Bézier-editorn  
Visar kontrollpunkterna för alla stödpunkter när du markerar en Bézierkurva.  
Om rutan inte är aktiverad visas bara kontrollpunkterna för en markerad punkt.  
Kontur för varje enskilt objekt  
%PRODUCTNAME visar konturerna för varje objekt med en streckad linje vid förflyttning.  
Då märker du redan vid förflyttningen om enskilda objekt kan kollidera med andra objekt vid målpositionen.  
Om rutan inte är aktiverad visar %PRODUCTNAME bara en begränsningsrektangel som omfattar alla markerade objekt.  
Raster  
Här kan du definiera raster för att skapa och flytta objekt.  
Om du har aktiverat stödrastret men vill flytta eller skapa enstaka objekt utan anpassning till stödrastret, håller du ner Kommando Ctrl -tangenten och sätter på så vis den här funktionen temporärt ur spel.  
Fäst  
Mot stödlinjer  
Med den här rutan justeras grafikobjektets kontur till närmaste stödlinje.  
Detta händer bara om muspekaren eller en av grafikobjektets konturlinjer befinner sig inom fästområdet.  
Ikonen finns på alternativlisten i ett öppet presentations - eller teckningsdokument.  
Mot sidmarginalerna  
Om du markerar den här rutan justeras grafikobjektets kontur till närmaste sidmarginal.  
Muspekaren eller en av grafikobjektets konturlinjer måste finnas inom fästområdet.  
Ikonen finns på alternativlisten när du har öppnat ett presentations - eller teckningsdokument.  
Mot objektram  
Om du markerar den här rutan justeras grafikobjektets kontur efter närmaste grafikobjekt.  
Muspekaren eller en av grafikobjektets konturlinjer måste finnas inom fästområdet.  
Ikonen finns på alternativlisten när du har öppnat ett presentations - eller teckningsdokument.  
Mot objektpunkter  
Grafikobjektets kontur justeras till närmaste grafikobjekts objektpunkter.  
Detta gäller bara då muspekaren eller en av grafikobjektets konturlinjer finns inom fästområdet.  
Ikonen finns på alternativlisten när du har öppnat ett presentations - eller teckningsdokument.  
Fästområde  
Med fästområdet definierar du avståndet mellan muspekaren och / eller objektkonturen.  
Detta avstånd måste underskridas för att %PRODUCTNAME Impress ska söka närmaste stödpunkt.  
Fästområdet definieras alltid i bildskärmspixel, det är oberoende av den valda skalan i vyn.  
Om du vill undvika för stora "hopp" när du skapar och placerar grafikobjekt, bör du inte öka fästområdets förvalda värde i för stora steg, bara från ca 5 till 10 pixel (bildpunkter).  
Anpassa till stödraster  
När objekt skapas och flyttas  
Grafikobjekt fixeras horisontellt, vertikalt eller diagonalt (45°) när de skapas eller flyttas.  
När du skapar en rektangel blir den därför en kvadrat och en ellips blir en cirkel.  
Om du tillfälligt vill sätta den här inställningen ur spel när du redigerar, håller du ner skifttangenten.  
Längre kantlängd  
Om du ritar upp en rektangel eller en ellips och sedan håller ned skifttangenten utan att släppa musknappen, skapas en kvadrat eller en cirkel med utgångspunkt från den längsta kanten.  
Om rutan Längre kantlängd inte är markerad, skapas kvadraten eller cirkeln med utgångspunkt från den kortare kanten.  
Vid rotation  
Grafikobjekt kan bara roteras runt den i textfältet angivna rotationsvinkeln.  
Om ett objekt ska roteras utöver den angivna vinkeln, håller Du ned Kommando Ctrl -tangenten under rotationen.  
När Du har uppnått önskad rotationsvinkel släpper Du tangenten.  
Punktreduktion  
I det här rotationsfältet definierar du vinkeln för punktreduktion.  
När du t.ex. redigerar polygoner kan du ha nytta av att reducera redigeringspunkterna i polygonen.  
Skriv ut  
Här väljer du vilka av teckningens eller presentationens element som ska skrivas ut.  
Tomma presentationsobjekt skrivs inte ut.  
Innehåll  
I det här området väljer du vilka delar av dokumentet som ska skrivas ut.  
Teckning  
Markera den här kryssrutan om sidans grafiska innehåll ska skrivas ut.  
Anteckningar  
Markera här om anteckningar ska skrivas ut.  
Flygblad  
Markera här om flygblad ska skrivas ut.  
Disposition  
Markera här om dispositionen ska skrivas ut.  
Utmatningskvalitet  
Standard  
Välj det här alternativet om du vill skriva ut med originalfärger.  
Gråskalor  
Välj det här alternativet om du vill skriva ut färger som gråskalor.  
Svartvitt  
Välj det här alternativet om du vill skriva ut dokumentet i svartvitt.  
Skriv ut  
I det här området väljer du de element som ska infogas i sidmarginalen då dokumentet skrivs ut.  
Du kan inte välja Sidnamn, Datum eller Tid när du har markerat Prospekt som sidalternativ.  
Sidnamn  
Markera detta alternativ om sidflikarnas namn ska skrivas ut.  
Datum  
Markera detta alternativ om det aktuella systemdatumet ska skrivas ut.  
Tid  
Markera detta alternativ om den aktuella systemtiden ska skrivas ut.  
Dolda sidor  
Markera här när du även vill skriva ut de sidor som du har dolt i presentationen.  
Sidalternativ  
I detta område anger Du ytterligare alternativ för hur utskriften av sidan ska se ut.  
Standard  
Markera detta alternativ om Du inte vill att sidornas storlek ska ändras vid utskrift.  
Anpassa till sidstorlek  
Välj det här alternativet så anpassas storleken på alla sidelement till sidstorleken vid utskrift.  
Sidor sida vid sida  
Välj det här alternativet när sidorna ska skrivas ut sida vid sida.  
Då måste du ha valt ett sidformat som är större än pappersformatet.  
Prospekt  
Välj det här alternativet när du vill skriva ut en broschyr.  
Du väljer om framsidan, baksidan eller båda sidorna ska skrivas ut.  
Bestäm först om du vill skriva på den ena eller båda sidorna.  
Om du vill skriva ut på en sida markerar du Framsida och Baksida och skriver sedan ut dem.  
Om du vill skriva på båda sidorna markerar du till att börja med bara Framsida och startar utskriften.  
Markera Baksida och fortsätt att skriva ut.  
Vik sidorna på mitten och prospektet är färdigt.  
Framsida  
Markera den här rutan om du vill skriva ut framsidorna i en broschyr.  
Baksida  
Markera den här rutan om du vill skriva ut baksidorna i en broschyr.  
Pappersfack från skrivarinställning  
Via detta alternativ anger du, för skrivare med flera pappersmagasin, om pappersmagasin ska väljas från skrivarens systeminställningar.  
Allmänt  
Här kan du göra allmänna inställningar.  
Du definierar t.ex. om textobjekt först ska markeras eller redigeras samt om en kopia ska skapas när du flyttar ett objekt.  
Textobjekt  
Tillåt snabbredigering  
Om den här rutan är markerad startar du textredigeringsläget när du klickar på en text i ett textobjekt.  
När ett presentations - eller teckningsdokument är öppet kan du också aktivera det här läget med hjälp av ikonen med samma namn på alternativlisten.  
Bara textområde kan markeras  
Det räcker inte att du klickar på ramen.  
I andra (ännu inte fyllda) områden kan du markera objekt som ligger under textramar.  
När ett presentations - eller teckningsdokument är öppet kan du också aktivera det här läget med hjälp av ikonen med samma namn på alternativlisten.  
Nytt dokument (bara för presentationer)  
Starta med AutoPiloten  
Aktivera den här rutan om du vill ha hjälp av AutoPiloten när du skapar en ny presentation via menyn Arkiv - Nytt - Presentation.  
Inställningar  
Här gör du fler inställningar.  
Använd cache för bakgrund  
Om du vill påskynda uppdateringen av bakgrunden kan du spara bakgrunden i cachen.  
Kopia vid förflyttning  
Markera den här rutan när du vill flytta (rotera, dimensionera) en kopia av originalet när du flyttar (roterar, dimensionerar) ett objekt genom att hålla ner Kommando Ctrl -tangenten.  
Originalet blir kvar på den ursprungliga platsen.  
Om du flyttar objekt utan att hålla ner tangenten flyttas bara originalet.  
Objekt alltid flyttbara  
När du redigerar ett teckningselement, t.ex. genom att rotera det, kan du samtidigt flytta teckningselementet.  
Om du vill stänga av den här dubbelfunktionen, avmarkerar du den här kryssrutan.  
Måttenhet  
Här väljer du måttenhet för presentationer.  
Tabulatoravstånd  
I det här rotationsfältet definierar du tabulatoravståndet.  
Sätt på cirkel: förvräng inte (bara för teckningar)  
Punkterna för tvådimensionella teckningselement och Bézierkurvor behåller sin justering till varandra även om du förvränger grafikobjektets perspektiv.  
Starta presentation (bara för presentationer)  
%PRODUCTNAME Impress startar presentationen antingen med den första sidan eller med den aktuella sidan.  
Alltid med aktuell sida  
Markera den här rutan när du vill att presentationen alltid ska starta med den aktuella sidan.  
Kompatibilitet (bara för presentationer)  
Här ställer du in kompatibiliteten till Microsoft PowerPoint-dokument.  
Addera alla styckeavstånd i det aktuella dokumentet  
Om den här rutan är markerad reagerar %PRODUCTNAME Impress precis som Microsoft PowerPoint när styckeavstånd beräknas.  
Microsoft PowerPoint adderar det övre och undre styckeavståndet. %PRODUCTNAME Impress använder bara det större av de båda.  
Skala (bara för teckningar)  
Teckningsskala  
Här väljer du teckningsskalan på linjalerna.  
Alternativ Teckning  
Här kan du göra olika globala inställningar för teckningsdokument.  
Bland annat definierar du vilket innehåll som ska visas på sidorna, vilken skala som ska gälla generellt, om, och i så fall hur, raster ska justeras och vilket innehåll som ska tas med vid utskrift.  
Skala  
Här anger du skalan för linjalerna.  
I programmet hanteras alltid sidstorleken i hundradels millimeter och här kan du ändra linjalenheternas förhållande till de interna enheterna.  
Efter Sidbredd och Sidhöjd visas sidstorleken som motsvarar det pappersformat som Du har valt.  
När Du ställer in en annan skala anpassas visningen av linjalerna till denna.  
Detta innebär att Du direkt kan kontrollera avstånden på papperet i de aktuella enheterna.  
Ange t ex skalan 1:50 när Du vill göra en planritning av vardagsrummet.  
På linjalerna ser Du nu att de inte längre motsvarar en yta på 29 gånger 21 centimeter, utan en yta på drygt 12 gånger 8 meter.  
Nu kan Du placera in och dimensionera objekten (t ex väggar, dörrar och fönster) med korrekta mått. (Eftersom bildskärmar för närvarnande inte är så stora att de kan visa flera metrar utan högst några dussin centimetrar kan det vara en bra idé att göra hela ritningen i centimeter i stället för meter.  
Detta ställer Du in direkt på linjalerna.)  
Skala  
I detta område ändrar Du skalan.  
När Du ändrar skalan anpassas storleken proportionellt i rotationsfälten Originalbredd och Originalhöjd.  
När Du ändrar något av de båda rotationsfälten anpassas på samma sätt inmatningen i fältet Skala så snart en passande skala uppnås.  
Skala  
I detta kombinationsfält väljer Du skala när Du vill ändra den proportionellt.  
Markera en av skalorna i listrutan eller ange själv en skala.  
När Du själv anger skalan kan Du t ex skriva 1:11 eller 7:1.  
Sidbredd  
Här visas sidbredden i den interna enheten 1 / 100 millimeter.  
Sidhöjd  
Här visas sidhöjden i den interna enheten 1 / 100 millimeter.  
Originalbredd  
I detta rotationsfält visas den beräknade nya originalbredden baserad på skalan.  
Du kan också ange ett eget värde om Du t ex vill ha olika skalor för bredd respektive höjd.  
Originalhöjd  
I detta rotationsfält visas den beräknade nya originalhöjden baserad på skalan.  
Du kan också ange ett eget värde om Du t ex vill ha olika skalor för bredd respektive höjd.  
Formel  
Här väljer du utskriftsformat och utskriftsalternativ för alla nya formeldokument.  
De här alternativen gäller om du vill skriva ut en formel direkt från %PRODUCTNAME Math.  
Du kan även öppna den här dialogrutan för den aktuella utskriften via kommandoknappen Fler i dialogrutan Skriv ut.  
Dina inställningar i dialogrutan Alternativ gäller permanent, medan inställningarna i dialogrutan "Skriv ut" bara gäller för det enstaka utskriftsjobbet.  
Inställningar  
Inställningar  
Här definierar du inställningar som ska gälla för alla dokument.  
Utskriftsalternativ  
Rubrikrad  
Markera den här rutan om rubriken som du angett då du sparade också ska skrivas ut.  
Formeltext  
Markera den här rutan om innehållet i fönstret Kommandon i den undre marginalen på utskriftssidan också ska skrivas ut.  
Ram  
Formelområdet på utskriften ramas in av en tunn heldragen linje.  
Utskriftsformat  
Här kan du definiera i vilken storlek formeln ska skrivas ut.  
Originalstorlek  
Formeln skrivs ut utan ändring i aktuell teckenstorlek.  
För större formler kan ibland en del av kommandotexten klippas av.  
Anpassa sida  
Formeln anpassas så att den fyller hela utskriftssidan.  
Den faktiska storleken bestäms av aktuellt pappersformat.  
Skalning  
Formeln förminskas eller förstoras med en viss procentfaktor vid utskrift.  
Ange önskad förstoringsfaktor direkt i rotationsfältet eller ställ in värdet med pilknapparna bredvid rotationsfältet.  
Övriga alternativ  
Ignorera ~ och 'vid radslutet  
Om du markerar den här kryssrutan tas de här platshållarna för blanksteg bort om de står vid ett radslut.  
Alternativ Diagram  
Här gör du allmänna förinställningar för dina diagram.  
Grundfärger  
Här definierar du dataseriernas färger.  
Inställningarna gäller bara för alla nya diagram.  
Diagramfärger  
Här visas alla inställda färger för dataserier.  
Markera en dataserie om du vill ändra dess färg.  
Välj en färg från färgtabellen som finns bredvid.  
Färgtabell  
Den här tabellen innehåller ersättning för diagramfärgerna i de markerade dataserierna.  
Om du exempelvis har markerat dataserie 6 och sedan klickar på färg Grön 8, ersätts dataseriens gamla färg med Grön 8.  
Namnet på den utvalda färgen visas under färgtabellen.  
Standard  
Med hjälp av den här kommandoknappen återställer du färginställningarna som gällde vid installationen.  
VBA-egenskaper  
Här gör du allmänna inställningar som gäller när du laddar och sparar Microsoft Office-dokument med VBA-kod.  
Microsoft Word 97 / 2000  
Här väljer du inställningarna för Microsoft Word 97 / 2000-dokument.  
Ladda Basic-kod för redigering  
Om den här rutan är markerad, laddas Basic-koden från Microsoft-dokumentet och sparas i särskild form som %PRODUCTNAME Basic-modul med dokumentet.  
Den noteras som kommentarer, inom parentes mellan Sub - och End Sub -kommandon.  
Du kan redigera koden.  
Om du sparar dokumentet i %PRODUCTNAME -format sparas Basic-koden med det.  
Om du sparar i ett annat format sparas inte Basic-koden från %PRODUCTNAME Basic-IDE:n.  
Spara original-Basic-kod igen  
Om den här rutan är aktiverad sparas Microsoft Basic-koden, som finns i dokumentet och är oförändrad, så länge i ett särskilt internt minne som dokumentet är laddat i %PRODUCTNAME.  
Om du sparar dokumentet i Microsoft-formatet sparas också Microsoft Basic oförändrat igen.  
Om du sparar i andra format än Microsoft-formatet går Microsoft Basic-koden förlorad.  
Om dokumentet innehåller Microsoft Basic-kod och du t.ex. sparar det i %PRODUCTNAME -format informerar dig ett varningsmeddelande om att Microsoft Basic-koden inte sparas.  
Om båda rutorna är aktiverade och du redigerar den kommenterade Basic-koden i %PRODUCTNAME Basic IDE:n, sparas original-Microsoft Basic-koden när du sparar i Microsoft-format.  
Ett meddelande informerar dig om detta.  
Tips: om du vill ta bort eventuella Microsoft Basic-makrovirus från Microsoft-dokumentet, avmarkerar du rutan Spara original-Basic-kod igen och sparar dokumentet i Microsoft-format.  
Dokumentet sparas då utan Microsoft Basic-kod.  
Microsoft Excel 97 / 2000  
Här väljer du inställningarna för Microsoft Excel 97 / 2000-dokument.  
Ladda Basic-kod för redigering  
Spara original-Basic-kod igen  
Microsoft PowerPoint 97 / 2000  
Här väljer du inställningarna för Microsoft PowerPoint 97 / 2000-dokument.  
Ladda Basic-kod för redigering  
Spara original-Basic-kod igen  
Microsoft Office  
Här gör du inställningar för import och export av Microsoft Office OLE-objekt.  
De här inställningarna gäller om det inte finns någon Microsoft OLE-server (t.ex. i UNIX) eller det inte finns någon %PRODUCTNAME OLE-server som kan redigera OLE-objekten.  
Listruta  
I listrutan finns poster för OLE-objektparen som kan omvandlas när de laddas i %PRODUCTNAME (L) och / eller när de sparas i ett Microsoft-format (S).  
Markera rutan i kolumnen [L] framför posten om ett Microsoft-OLE-objekt ska omvandlas till det nämnda %PRODUCTNAME -OLE-objektet när ett Microsoft-dokument laddas i %PRODUCTNAME.  
Markera rutan i kolumnen [S] framför posten om ett %PRODUCTNAME -OLE-objekt ska omvandlas till det nämnda Microsoft-OLE-objektet när ett dokument sparas i ett Microsoft-filformat.  
Språk  
Här väljer du bl.a. standardspråken för dokumenten.  
Språk för  
Språkvariant  
Här väljer du språkvarianten (locale) av landsinställningen.  
Den påverkar inställningar för tal, valuta och måttenheter.  
Posten "standard" står för språkvarianten som har valts för operativsystemet.  
En ändring i den här rutan träder i kraft direkt.  
Men talformat som har formaterats som "standard" ändras först när dokumentet laddas om på nytt.  
Standardvaluta  
Här väljer du standardvalutan som t.ex. används för valutaformatet och för valutafälten.  
Om du byter språkvariant byts även standardvalutan automatiskt.  
Posten "standard" står för valutaformatet som har tilldelats den valda språkvarianten.  
En ändring i den här rutan överförs till alla öppnade dokument och leder till en motsvarande ändring i dialogrutorna och ikonerna som styr valutaformatet.  
Standardspråk för dokument  
Här väljer du språken t.ex. för rättstavningskontroll, synonymordlista och avstavning.  
Rättstavningskontroll för det valda språket fungerar bara om du har installerat motsvarande språkmodul.  
Västligt  
Här definierar du vilket språk som ska användas för rättstavningskontrollen i västliga alfabet.  
Asiatiskt  
Här definierar du vilket språk som ska användas för rättstavningskontrollen i asiatiska alfabet.  
Bara för det aktuella dokumentet  
Markera den här rutan om inställningarna i det här området bara ska gälla för det aktuella dokumentet.  
Stöd för asiatiska språk  
%PRODUCTNAME stöder specialfunktionerna för asiatiska språk med många inställningar i många dialogrutor.  
Om du aldrig skriver på kinesiska, japanska eller koreanska kan du ta bort stödet från programgränssnittet.  
Aktiverat  
Markera den här rutan om du även vill göra inställningar för asiatiska språk i motsvarande dialogrutan.  
Alternativ språkinställningar  
Här bestämmer du egenskaperna för språk.  
Sökalternativ för japanska och Asiatisk layout ser du bara om du har aktiverat Stöd för asiatiska språk under Språk och har öppnat Alternativ-dialogrutan på nytt.  
Asiatisk layout  
Här väljer du typografiska förinställningar för asiatiska texter.  
Kerning  
Här gör du förinställningar för minskning av mellanrum mellan enskilda tecken (kerning).  
Bara västliga tecken  
Om du väljer det här alternativet används kerning bara för västlig text.  
Västliga tecken och asiatisk interpunktion  
Om du väljer det här alternativet används kerning för västlig text och asiatisk interpunktion.  
Teckenavstånd  
Här gör du förinställningar för teckenavståndet i asiatiska texter, cellinnehåll och ritobjekt.  
Ingen kompression  
Om du väljer det här alternativet sker ingen kompression.  
Komprimera bara interpunktion  
Om du väljer det här alternativet komprimeras bara interpunktionen.  
Komprimera interpunktion och japansk Kana  
Om du väljer det här alternativet komprimeras interpunktionen och japansk Kana.  
Start - och sluttecken  
Här gör du förinställningar för start - och sluttecken.  
I dialogrutan Format under fliken Asiatisk typografi definierar du för stycket eller för styckeformatmallen om listan med förbjudna tecken i början och slutet av raden används för ett stycke.  
Språk  
Här väljer du språket.  
De språk vars lingvistik är installerade i ditt %PRODUCTNAME har en grön markering.  
Standard  
Markera den här rutan om språkvalet ska gälla som standard.  
Inte i början av rad:  
Här matar du in de tecken som inte får stå ensamma i början av en rad.  
Om ett av de här tecknen skulle hamna i början av raden vid en brytning flyttas det automatiskt till slutet av föregående rad.  
Ett utropstecken efter det sista ordet i en mening kommer till exempel aldrig att stå i början av en rad om du matar in det här.  
Inte i slutet av rad:  
Här matar du in de tecken som inte får stå ensamma i slutet av en rad.  
Om ett av de här tecknen skulle hamna i slutet av raden vid en brytning flyttas det automatiskt till början av nästa rad.  
Ett valutatecken som står framför valutabeloppet kommer till exempel aldrig att stå i slutet av en rad om du matar in det här.  
Sökalternativ för japanska  
Här väljer du sökalternativen för japanska.  
Behandla likvärdigt  
Här väljer du alternativet som ska behandlas likvärdigt i en sökning.  
Ignorera  
Här väljer du tecknet som ska ignoreras.  
Alternativ Datakällor  
Här gör du allmänna förinställningar för datakällorna i %PRODUCTNAME.  
Förbindelser  
Här definierar du hur poolningen av datakällor ska göras.  
Att skapa en anslutning till en datakälla kostar resurser och tid.  
Därför kan du ställa in här att anslutningarna som inte längre används inte raderas direkt utan hålls kvar en stund.  
Om en ny anslutning behövs under den här tiden kan anslutningen som har blivit ledig användas till det.  
Poolning av kopplingar  
Om den här rutan är markerad sker poolning av de anslutningar som du väljer.  
Om den här rutan inte är markerad sker ingen poolning av någon anslutning.  
Kända drivrutiner i %PRODUCTNAME  
Här ser du listan med drivrutiner och kopplingsdata som du har definierat.  
Poolning av kopplingar för den här drivrutinen  
Välj en drivrutin i listan och markera den här rutan för att poolning ska göras för den.  
Timeout (sekunder)  
Om poolning görs för en anslutning kan du välja hur länge anslutningen ska hållas kvar i sekunder.  
Tiden kan ligga mellan 30 och 600 sekunder.  
Så hittar du den här funktionen...  
Menyn Redigera  
Menyn Redigera - Sidhuvud och sidfot...  
Menyn Redigera - Sidhuvud och sidfot... - fliken Sidhuvud / sidfot  
Menyn Redigera - Ifyllning  
Menyn Redigera - Ifyllning - NedÃ¥t  
Menyn Redigera - Ifyllning - HÃ¶ger  
Menyn Redigera - Ifyllning - UppÃ¥t  
Menyn Redigera - Ifyllning - VÃ¤nster  
Menyn Redigera - Ifyllning - Tabell...  
Menyn Redigera - Ifyllning - Serie...  
Menyn Redigera - Radera innehåll...  
Tangenten Delete  
Menyn Redigera - Radera celler...  
Menyn Redigera - Radera tabell...  
Snabbmenyn på tabellflikarna  
Menyn Redigera - Kopiera / Flytta tabell...  
Snabbmenyn på tabellflikarna  
Menyn Redigera - Radera manuell brytning  
Menyn Redigera - Radera manuell brytning - Radbrytning  
Menyn Redigera - Radera manuell brytning - Kolumnbrytning  
Menyn Visa  
Menyn Visa - Kolumn - / radhuvuden  
Menyn Visa - FramhÃ¤v vÃ¤rden  
Menyn Visa - Symbollister - Formellist  
Menyn Visa - FÃ¶rhandsvisning av sidbrytningar  
Menyn Infoga  
Menyn Infoga - Manuell brytning  
Menyn Infoga - Manuell brytning - Radbrytning  
Menyn Infoga - Manuell brytning - Kolumnbrytning  
Menyn Infoga - Celler...  
Ikon på utrullningslisten Infoga celler på verktygslisten:  
Infoga celler  
Infoga celler, nedåt  
Infoga celler, till höger  
Infoga rader  
Infoga kolumner  
Menyn Infoga - Rader  
Menyn Infoga - Kolumner  
Menyn Infoga - Tabell...  
Menyn Infoga - Funktion...  
Tangentkombinationen Kommando Ctrl +F2  
Ikon på formellisten:  
Funktionsautopilot  
Funktionsautopilot - kategori Databas  
Funktionsautopilot - kategori Datum&Tid  
Funktionsautopilot - kategori Finans  
Funktionsautopilot - kategori Information  
Funktionsautopilot - kategori Logisk  
Funktionsautopilot - kategori Matematik  
Funktionsautopilot - kategori Matris  
Funktionsautopilot - kategori Statistik  
Funktionsautopilot - kategori Text  
Funktionsautopilot - kategori Tabell  
Funktionsautopilot - kategori Add-In  
Funktionsautopilot - kategori Add-in  
Menyn Infoga - Funktionslista  
Menyn Infoga - Namn  
Menyn Infoga - Externa data...  
Menyn Infoga - Namn - Definiera...  
Tangentkombinationen Kommando Ctrl +F3  
Menyn Infoga - Namn - Klistra in...  
Menyn Infoga - Namn - Ã–verta...  
Menyn Infoga - Namn - Etiketter...  
Menyn Format  
Menyn Format - Cell...  
Menyn Format - Cell... - fliken Cellskydd  
Menyn Format - Rad  
Menyn Format - Rad - Optimal hÃ¶jd...  
Menyn Format - Rad - Dölj  
Menyn Format - Kolumn - Dölj  
Menyn Format - Tabell - Dölj  
Menyn Format - Rad - Visa  
Menyn Format - Kolumn - Visa  
Menyn Format - Kolumn  
Menyn Format - Kolumn - Optimal bredd...  
Ikon på objektlisten:  
Dubbelklicka på den högra kolumnavgränsaren i kolumnhuvudena  
Menyn Format - Tabell  
Menyn Format - Tabell - Byt namn...  
Menyn Format - Tabell - Visa...  
Menyn Format - Sammanfoga celler  
Menyn Format - Sammanfoga celler - Definiera  
Menyn Format - Sammanfoga celler - UpphÃ¤v  
Menyn Format - Sida...  
Dubbelklicka på fältet på statuslisten  
Ikon på förhandsgranskningslisten:  
Sidformat  
Menyn Format - Sida... - fliken Tabell  
Menyn Format - UtskriftsomrÃ¥den  
Menyn Format - UtskriftsomrÃ¥den - Definiera  
Menyn Format - UtskriftsomrÃ¥den - LÃ¤gg till  
Menyn Format - UtskriftsomrÃ¥den - UpphÃ¤v  
Menyn Format - UtskriftsomrÃ¥den - Redigera  
Menyn Format - Mallkatalog...  
Tangentkombinationen Kommando Ctrl +Y  
Menyn Format - AutoFormat...  
Ikon på verktygslisten:  
AutoFormat  
Menyn Format - Villkorlig formatering...  
Menyn Verktyg  
Menyn Verktyg - Detektiv  
Menyn Verktyg - Detektiv - Spåra föregångare  
Tangentkombinationen Ctrl+F5  
Menyn Verktyg - Avstavning  
Menyn Verktyg - Detektiv - Ta bort spÃ¥r till fÃ¶regÃ¥ngare  
Menyn Verktyg - Detektiv - Spår till efterträdaren  
Tangentkombinationen Skift+F5  
Menyn Verktyg - Detektiv - Ta bort spÃ¥r till eftertrÃ¤dare  
Menyn Verktyg - Detektiv - Ta bort alla spÃ¥r  
Menyn Verktyg - Detektiv - SpÃ¥r till fel  
Menyn Verktyg - Detektiv - FyllningslÃ¤ge  
Menyn Verktyg - Detektiv - Ringa in ogiltiga data  
Menyn Verktyg - Detektiv - Uppdatera spÃ¥r  
Menyn Verktyg - Detektiv - Uppdatera automatiskt  
Menyn Verktyg - MÃ¥lvÃ¤rdessÃ¶kning...  
Menyn Verktyg - Scenarion...  
Menyn Verktyg - Skydda dokument  
Menyn Verktyg - Skydda dokument - Tabell...  
Menyn Verktyg - Skydda dokument - Dokument...  
Menyn Verktyg - CellinnehÃ¥ll  
Menyn Verktyg - Cellinnehåll - Beräkna på nytt  
Tangenten F9  
Menyn Verktyg - CellinnehÃ¥ll - Automatisk berÃ¤kning  
Menyn Verktyg - CellinnehÃ¥ll - AutoInmatning  
Menyn Fönster  
Menyn FÃ¶nster - Dela  
Menyn FÃ¶nster - Fixera  
Menyn Data  
Menyn Data - Definiera omrÃ¥de...  
Menyn Data - VÃ¤lj omrÃ¥de...  
Menyn Data - Sortera...  
Menyn Data - Sortera - fliken Sorteringskriterier  
Ikoner på verktygslisten:  
Sortera stigande  
Sortera fallande  
Menyn Data - Sortera - fliken Alternativ  
Menyn Data - Filter  
Menyn Data - Filter - AutoFilter  
Ikon på verktygslisten och på databaslisten:  
Automatiskt filter  
Menyn Data - Filter - Specialfilter...  
Menyn Data - Filter - Standardfilter... - kommandoknappen Fler  
Menyn Data - Filter - Specialfilter... - kommandoknappen Fler  
Menyn Data - Filter - Ta bort filter  
Databaslisten - ikonen Ta bort filter / sortering  
Ta bort filter / sortering  
Menyn Data - Filter - DÃ¶lj AutoFilter  
Menyn Data - Delresultat...  
Menyn Data - Delresultat... - flikarna Grupp 1, 2, 3  
Menyn Data - Delresultat... - fliken Alternativ  
Menyn Data - Validitet...  
Menyn Data - Validitet - fliken Kriterier  
Menyn Data - Validitet... - fliken InmatningshjÃ¤lp  
Menyn Data - Validitet... - fliken Felmeddelande  
Menyn Data - Multipla operationer...  
Menyn Data - Konsolidera...  
Menyn Data - Disposition  
Menyn Data - Disposition - DÃ¶lj detalj  
Menyn Data - Disposition - Visa detalj  
Menyn Data - Disposition - Gruppering...  
Tangenten F12  
Ikon på verktygslisten:  
Infoga gruppering  
Menyn Data - Disposition - Upphäv gruppering...  
Tangentkombinationen Kommando Ctrl +F12  
Ikon på verktygslisten:  
Ta bort gruppering  
Menyn Data - Disposition - AutoDisposition  
Menyn Data - Disposition - Ta bort  
Menyn Data - Datapilot  
Menyn Data - Datapilot - Starta...  
Menyn Data - Datapilot - Starta... - Välj ut källa - alternativet Datakälla som är registrerad i %PRODUCTNAME  
Menyn Data - Datapilot - Starta... - Välj ut källa - alternativet Aktuell markering  
Menyn Data - Datapilot - Starta... - Välj ut källa - alternativet Datakälla som är registrerad i %PRODUCTNAME - VÃ¤lj ut datakÃ¤lla  
Menyn Data - Datapilot - Uppdatera  
Menyn Data - Datapilot - Radera  
Menyn Data - Uppdatera omrÃ¥de...  
Navigator  
Här kan du visa och dölja Navigator.  
Navigator är ett förankringsbart fönster.  
Om du vill att Navigator ska visas på bildskärmen, väljer du Redigera - Navigator när ett dokument är öppet, klickar på ikonen på funktionslisten eller trycker på F5.  
Du kan flytta Navigator-fönstret genom att placera muspekaren på titellisten, hålla ner musknappen och dra fönstret.  
Om Navigator-fönstret ska förankras vid fönsterkanten när du flyttar det, håller du ner Kommando Ctrl -tangenten.  
Kolumn  
I detta rotationsfält kan du ange en kolumnbokstav.  
Den stannar dock kvar på samma rad.  
Rad  
I det här rotationsfält et kan du ange ett radnummer.  
Den stannar dock kvar i samma kolumn.  
Dataområde  
Via detta alternativ markerar %PRODUCTNAME Calc det aktuella dataområdet, beroende på cellmarkörens position.  
Dataområde  
Början  
Via den här ikonen kommer du till början av det aktuella dataområdet som du kan framhäva med kommandoknappen Dataområde.  
Början  
Slut  
Via den här ikonen kommer du till slutet av det aktuella dataområdet som du kan framhäva med kommandoknappen Dataområde.  
Slut  
Växla  
Med denna ikon växlar du innehållsvy.  
Det element som är markerat i Navigator görs till ursprung för visningen i Navigator och sedan visas bara detta element och dess underordnade element.  
Om du klickar på ikonen på nytt visas vyn med alla element igen.  
Växla  
Innehåll  
Här kan du visa och dölja visningen av innehållet.  
Innehåll  
Scenarion  
Här visas de definierade namnen på scenarion.  
Du kan använda ett scenario genom att dubbelklicka på dess namn.  
I tabellen visas sedan resultatet av ditt val.  
Ytterligare information får du via menyn Verktyg - Scenarion.  
Scenarion  
Draläge  
Med den här ikonen väljer du draläget.  
Om du klickar på ikonen och håller ner musknappen visas en undermeny, där du kan välja mellan följande lägen:  
Draläge  
Infoga som hyperlänk  
Draläget hyperlänk infogar en hyperlänk vid dra-och-släpp från Navigator.  
Infoga som länk  
Draläget länk infogar en länk via dra-och-släpp från Navigator.  
Infoga som kopia  
Draläget kopia infogar en kopia via dra-och-släpp från Navigator.  
Existerande objekt  
I det här området visas en lista över alla objekt som finns i dokumentet.  
Dokumentlista  
I det här kombinationsfältet visas namnen på de laddade dokumenten.  
Om du vill växla till ett annat laddat dokument i Navigator, klickar du på dokumentnamnet.  
Efter varje dokumentnamn visas inom parentes om dokumentet är aktivt eller inaktivt.  
Det aktiva dokumentet väljer du på menyn Fönster.  
Sidhuvuden och sidfötter  
Med det här kommandot kan du definiera och formatera sidhuvuden och sidfötter.  
Den här dialogrutan innehåller flikar där du definierar sidhuvuden och sidfötter.  
Om du har angett att innehållet på höger - och vänstersidor inte ska vara detsamma i dialogrutan Sidformatmall, visas skilda flikar för dokumentets vänstersidor och högersidor.  
Sidhuvud / sidfot  
Här kan du definiera eller formatera en sidhuvud / sidfot för en sidformatmall.  
Vänster område  
Här kan du ange en text som ska visas till vänster i sidhuvudet / sidfoten.  
Mittområde  
Här kan du ange en text som ska visas centrerat i sidhuvudet / sidfoten.  
Höger område  
Här kan du ange en text som ska visas till höger i sidhuvudet / sidfoten.  
Textattribut  
Här bestämmer du med vilka attribut den markerade texten, eller den nya text som skrivs in, ska formateras.  
Dialogrutan som öppnas innehåller flikarna Teckensnitt, Teckeneffekt och Teckenposition.  
Textattribut  
Filnamn  
Här kan du infoga en platshållare för filnamnet i det aktuella sidhuvuds - / sidfotsområdet.  
Detta gör det möjligt att visa filnamnet i det aktuella dokumentets sidhuvud / sidfot.  
Om du klickar snabbt infogas rubriken.  
Om du klickar litet längre visas en undermeny där du kan ange om rubrik, filnamn eller sökväg / filnamn ska infogas.  
Om du ännu inte gett dokumentet en rubrik (under Arkiv - Egenskaper) visas filnamnet istället för rubriken.  
Filnamn  
Tabellnamn  
Här kan du infoga en platshållare för tabellnamnet i det aktuella sidhuvuds - / sidfotsområdet.  
Detta gör det möjligt att visa tabellnamnet i sidhuvudet / sidfoten i det aktuella dokumentet.  
Tabellnamn  
Sida  
Här kan du infoga en platshållare för aktuellt sidnummer i det valda sidhuvuds - / sidfotsområdet.  
På så vis får du en löpande sidnumrering i dokumentet.  
Sida  
Sidor  
Här kan du infoga en platshållare för totalt antal sidor i det aktuella sidhuvuds - / sidfotsområdet.  
Totalt antal sidor i dokumentet visas i sidhuvuds - / sidfotsområdet.  
Sidor  
Datum  
Här kan du infoga en platshållare för aktuellt datum i det aktuella sidhuvuds - / sidfotsområdet.  
Aktuellt datum visas i sidhuvuds - / sidfotsområdet på alla sidor i dokumentet.  
Datum  
Klockslag  
Här kan du infoga en platshållare för aktuellt klockslag i det aktuella sidhuvuds - / sidfotsområdet.  
Aktuellt klockslag visas i sidhuvuds - / sidfotsområdet på alla sidor i dokumentet.  
Klockslag  
Fyll  
Med det här kommandot kan du fylla celler med innehåll automatiskt.  
Förutom att du kan använda kommandona på undermenyerna har du även en annan möjlighet att fylla i celler med hjälp av snabbmenyn i %PRODUCTNAME Calc.  
Tabell...  
Serie...  
Så här fyller du i celler via snabbmenyn:  
Öppna snabbmenyn i cellen och välj Urvalslista.  
Alla textposter i den aktuella kolumnen visas i en listruta.  
Textposterna är sorterade i bokstavsordning och eventuella dubbletter visas bara som en post i listan.  
Klicka på den post i listan som du vill överföra till den aktuella cellen.  
Nedåt  
Här kan du fylla ett markerat område som omfattar minst två rader med innehållet i den översta cellen i området.  
Om du bara har markerat en kolumn i ett område, kopieras innehållet i den översta cellen till alla andra celler i det markerade området.  
Om du har markerat flera kolumner, kopieras den översta cellen i varje kolumn till cellerna nedanför.  
Höger  
Här kan du fylla ett markerat område som omfattar minst två kolumner med innehållet i cellen som står längst till vänster.  
Om du bara har markerat en rad i ett område, kopieras innehållet i cellen längst till vänster till alla andra celler i det markerade området.  
Om du har markerat flera rader, kopieras cellen längst till vänster i varje rad till cellerna till höger om den.  
Uppåt  
Här kan du fylla ett markerat område, som omfattar minst två rader, med innehållet i den nedersta cellen.  
Om du har markerat ett område med bara en kolumn, kopieras innehållet i den nedersta cellen till alla andra celler i det markerade området.  
Om du har markerat flera kolumner kopieras den nedersta cellen i varje kolumn till cellerna ovanför.  
Vänster  
Här kan du fylla ett markerat område, som omfattar minst två kolumner, med innehållet i cellen längst till höger.  
Om ett område med bara en cell är markerat så kopieras innehållet i cellen längst till höger till alla andra celler inom det markerade området.  
Om flera rader är markerade kopieras innehållet i cellen längst till höger på varje rad till cellerna till vänster.  
Fyll tabeller  
Här väljer du bland olika alternativ för överföring av hela tabeller eller delområden i ett tabelldokument.  
Till skillnad från när du kopierar områden via urklippet kan du filtrera bort viss information och använda räkneoperationer på värdena.  
Det här kommandot är bara aktivt om dokumentet innehåller minst två markerade tabeller.  
Då måste du klicka på tabellfliken och samtidigt hålla ner Kommando Ctrl -tangenten eller skifttangenten, så att fliken framhävs mot ljus bakgrund.  
Så här fyller du en tabell  
Markera en hel tabell (klicka på rutan uppe till vänster i hörnet) eller tabellområdet i arbetsbladet som du vill överföra.  
Markera därefter tabellfliken till den aktuella tabellen där du vill infoga innehållet.  
Välj sedan Redigera - Fyll - Tabell....  
Om du vill knyta räkneoperationer till värdena måste du förstås ha markerat Siffror (eller Klistra in allt) i området Urval.  
Välj Räkneoperation vid behov.  
Klicka sedan på OK.  
Den här dialogrutan motsvarar innehållsmässigt tabelldokumentsdelen i dialogrutan Klistra in innehåll, där det finns ytterligare information.  
Fyll serier  
Med alternativen i den här dialogrutan kan du generera serier automatiskt.  
Du kan ange riktning, inkrement, tidsenhet och serietyp.  
Innan du fyller en serie måste det cellområde som ska fyllas vara markerat.  
I så fall ska du använda alternativet Serie med AutoFyll.  
Riktning  
I det här området kan du ange i vilken riktning serien ska skapas.  
Nedåt  
Här skapar du inom det markerade cellområdet en serie nedåt i kolumnen med angivet inkrement fram till maxvärdet.  
Höger  
Här skapar du inom det markerade cellområdet en serie som går från vänster till höger och med angivet inkrement fram till maxvärdet.  
Uppåt  
Här skapar du inom det markerade cellområdet uppåt i kolumnen en serie med angivet inkrement fram till maxvärdet.  
Vänster  
Här skapar du inom det markerade cellområdet en serie som går från höger till vänster och med angivet inkrement fram till maxvärdet.  
Serietyp  
I det här området kan du välja mellan serietyperna Aritmetisk, Geometrisk, Datum och AutoFyll.  
Aritmetisk  
Om det här alternativet är markerat, skapas en aritmetisk talserie på basis av angivet inkrement och maxvärdet.  
Geometrisk  
Om det här alternativet är markerat, skapas en geometrisk talserie på basis av angivet inkrement och maxvärdet.  
Datum  
Om det här alternativet är markerat, skapas en datumserie på basis av angivet inkrement och maxdatum.  
AutoFyll  
Du kan skapa en serie direkt i tabellen genom att använda AutoFyll.  
Den baseras då på användardefinierade listor.  
Om du t.ex. anger jan i den första cellen, fylls övriga celler automatiskt i enligt den lista som du har definierat under Verktyg - Alternativ - Tabelldokument - Sorteringslistor.  
AutoFyll fortsätter värdeserier enligt befintligt mönster.  
Exempelvis fortsätts serien 1, 3, 5 med 7, 9, 11, 13 osv.  
Serien 1, 3, 6 däremot fortsätts med 2, 4, 7, 3, 5, 8, 4, 6, 9 osv.  
Datum - och klockslagsserier fortsätts på motsvarande sätt; efter 1997-01-01 och 1997-01-15 räknas alltså vidare med 14-dagarsintervall.  
Tidsenhet  
I det här området kan du välja tidsenheterna Dag, Veckodag, Månad och År.  
Det här området är bara aktivt om du har markerat alternativet Datum i området Serietyp.  
Dag  
Om du har aktiverat Datum som serietyp, kan du skapa en serie med sjudagarsräkning.  
Veckodag  
Här kan du skapa en serie med femdagarsräkning, d.v.s. utan att veckosluten inkluderas.  
Månad  
Om serietypen Datum är aktiverad, kan du skapa en serie med månadsnamn eller månadsförkortningar.  
År  
Om serietypen Datum är aktiverad, kan du skapa en serie med årtal.  
Startvärde  
Här anger du startvärdet för serien som ska skapas.  
Det kan anges som tal, datum eller klockslag.  
Maxvärde  
Här anger du slutvärdet för den serie som ska skapas.  
Det kan anges som tal, datum eller klockslag.  
Inkrement  
Med termen "inkrement" menas det tal med vilket en storhet ökar.  
Ange i fältet värdet med vilket serien som du skapar ska ökas för varje steg, med hänsyn tagen till den valda serietypen.  
Du kan bara ange ett värde om du har valt serietypen Aritmetisk, Geometrisk eller Datum.  
Radera innehåll  
Här anger du vilket innehåll som ska raderas i en cell eller ett cellområde.  
Det är bara innehållet i markerade celler eller den aktuella cellen som raderas.  
Om du har markerat flera tabeller är det bara i den aktuella tabellen som raderingen sker.  
Den här dialogrutan kan du även öppna genom att trycka på Delete-tangenten på tangentbordet om cellmarkören samtidigt är aktiverad i tabellen.  
Formaten finns däremot kvar.  
Med ikonen Klipp ut på funktionslisten raderar du både innehåll och format utan att dialogrutan öppnas.  
Urval  
I det här området kan du välja vilket innehåll som ska raderas.  
Radera allt  
Om du markerar den här rutan raderas allt innehåll från det markerade cellområdet.  
Strängar  
Om du markerar den här rutan raderas bara strängar.  
Format och formler blir kvar.  
Siffror  
Om du markerar den här rutan raderas bara siffror.  
Format och formler blir kvar.  
Datum och tid  
Om du markerar den här rutan raderas bara datum och klockslag.  
Format, text, tal och formler blir kvar.  
Formler  
Om du markerar den här rutan raderas bara formler.  
Text, tal, format, datum och klockslag blir kvar.  
Anteckningar  
Om du markerar den här rutan raderas bara anteckningar som du har lagt till i cellerna.  
Alla andra element blir kvar.  
Format  
Om du markerar den här rutan raderas bara cellernas formatattribut.  
Allt innehåll finns kvar.  
Objekt  
Allt innehåll i cellerna finns kvar.  
Radera celler  
Här raderar du markerade celler, rader eller kolumner i sin helhet.  
Om du öppnar dialogrutan på nytt är det här alternativet markerat.  
Urval  
I det här området kan du välja hur tabellen ska se ut när cellerna har raderats.  
Flytta celler uppåt  
Klicka här om du vill att de celler som ligger under cellerna som ska raderas ska flyttas uppåt efter raderingen.  
Flytta celler åt vänster  
Klicka här om du vill att de celler som ligger till höger om cellerna som ska raderas ska flyttas åt vänster efter en radering.  
Radera hela rader  
Här kan du fullständigt radera en hel rad, där du markerat minst en cell, från tabellen.  
Radera hela kolumner  
Klicka här om du vill radera en hel kolumn, där du markerat minst en cell, från tabellen.  
Radera tabell  
Här kan du, efter en säkerhetskontroll, radera den aktuella tabellen.  
Observera att du inte kan radera en tabell om ändringar i dokumentet registreras, d.v.s. om menykommandot Redigera - Ändringar - Registrera är aktivt.  
Ja  
Om du vill radera den aktuella tabellen bekräftar du det genom att klicka på den här kommandoknappen.  
Nej  
Om du inte vill radera den aktuella tabellen bekräftar du det genom att klicka på den här kommandoknappen.  
Kopiera / Flytta tabell  
I den här dialogrutan kan du bestämma om du vill flytta eller kopiera den aktuella tabellen.  
Du kan flytta respektive kopiera tabellen inom dokumentet eller till ett annat dokument.  
Till dokument  
I det här kombinationsfältet kan du välja ett filnamn för ett öppnat dokument till vilket den aktuella tabellen ska flyttas eller kopieras.  
Välj alternativet - nytt dokument - om du vill skapa ett nytt dokument för den tabell som ska flyttas respektive kopieras.  
Infoga framför  
Välj namnet på en tabell framför vilken den aktuella tabellen ska flyttas resp. kopieras.  
Du kan också välja alternativet - flytta till slutet - om den aktuella tabellen ska flyttas till slutet.  
Kopiera  
Med det här alternativet bestämmer du om en tabell ska flyttas eller kopieras.  
Om du har markerat alternativet, så kopieras den aktuella tabellen.  
Standardinställningen är att tabeller flyttas.  
Radera manuell brytning  
Med det här kommandot öppnar du en undermeny, där du kan välja vilken typ av manuell radbrytning som ska raderas: radbrytning eller kolumnbrytning.  
Radbrytning  
Här kan du ta bort en manuell radbrytning direkt ovanför den aktuella cellen.  
Välj det här kommandot.  
Den manuella radbrytningen raderas.  
Kolumnbrytning  
Här kan du ta bort en manuell kolumnbrytning omedelbart till vänster om den aktuella cellen.  
Placera cellmarkören i en cell omedelbart till höger om kolumnbrytningen som är markerad med ett vertikalt streck.  
Den manuella kolumnbrytningen raderas.  
Kolumn - / radhuvuden  
Om du har markerat det här menyalternativet, visas tabellerna med kolumn - och radhuvuden.  
Om du vill dölja kolumn - och radhuvudena, avmarkerar du menyalternativet.  
Du kan också ställa in visningen av kolumn - och radhuvuden under Verktyg - Alternativ - Tabelldokument - Vy.  
Framhäv värden  
Om du aktiverar den här menyposten framhävs värdena i en tabell med färg.  
Om du vill stänga av färgsättningen, avmarkerar du menyposten.  
Textceller formateras med svart färg, celler som innehåller tal är blå och andra celler (formler, logiska värden, datum etc) är gröna.  
När detta kommando är aktivt visas inte de färger som har angetts i dokumentet.  
Färgerna finns dock kvar och visas igen när Du avmarkerar kommandot.  
Formellist  
Om det här menyalternativet är markerat, visas formellisten.  
Den är till för inmatning och redigering av formler och är det viktigaste verktyget när Du arbetar med tabelldokument.  
Du kan dölja formellisten genom att ta bort markeringen framför menyalternativet (klicka på det).  
Även om formellisten inte syns kan du redigera innehållet i den aktuella cellen om du går över till redigeringsläget genom att trycka på funktionstangenten F2.  
Redigera innehållet eller skriv över det (du behöver inte markera det) med ett nytt innehåll.  
Du ignorerar ändringen med Esc-tangenten.  
I så fall lämnar du även redigeringsläget.  
Förhandsvisning av sidbrytningar  
När du har markerat den här menyposten visas sidbrytningarna inne i tabellen.  
I förhandsvisningsläget för sidbrytningar gäller följande inställningar:  
Visningsskalan ställs in på 60%.  
Den del av tabellen som inte skrivs ut förses med en grå bakgrund.  
I mitten av varje utskriftssida visas sidnumret.  
Sidorna räknas inom tabellen från sida 1.  
Utskriftsområden och sidbrytningar visas med blå linjer.  
Mörkblå linjer markerar "automatiska" utskriftsområden och sidbrytningar.  
De markerar alltså den använda delen av tabellen om Du inte har definierat något utskriftsområde, och de markerar automatiskt insatta sidbrytningar.  
Manuellt definierade utskriftsområden och sidbrytningar visas i ljusblå färg.  
Du kan flytta de visade utskriftsområdena och sidbrytningarna med musen.  
När Du förminskar ett utskriftsområde så mycket att det inte finns något kvar, upphävs utskriftsområdet.  
Om det inte längre finns något utskriftsområde definierat för någon av tabellerna i dokumentet, så omfattar utskriften åter den del av tabellerna där det finns data.  
Om du flyttar en automatisk sidbrytning, så infogas en manuell brytning vid slutpositionen.  
Om Du flyttar en automatisk sidbrytning mot höger eller nedåt, så förminskas vid behov skalan så mycket att området mellan den flyttade och den tidigare brytningen ryms på en sida.  
Den ursprungliga brytningen förvandlas till en manuell brytning.  
Om Du flyttar en manuell sidbrytning utanför utskriftsområdet raderas den.  
På sidbrytningsförhandsvisningens snabbmeny hittar Du de viktigaste funktionerna för att redigera sidindelningen, bl a följande:  
Radera alla manuella brytningar  
Raderar alla manuella brytningar i den aktuella tabellen.  
Lägg till utskriftsområde  
Lägger till de markerade cellerna i tabellens befintliga utskriftsområden.  
Manuell brytning  
Här väljer du vilken typ av sidbrytning som ska infogas.  
En horisontell sidbrytning kan infogas ovanför den aktuella cellen, en vertikal sidbrytning till vänster om den aktuella cellen.  
Du tar bort en manuell brytning via menykommandot Redigera - Radera manuell brytning.  
Radbrytning  
Med det här kommandot infogar du en radbrytning (horisontell sidbrytning) ovanför den markerade cellen.  
Du känner igen en manuell radbrytning på den mörkblå horisontella linjen i tabellen.  
Kolumnbrytning  
Med det här kommandot infogar du en kolumnbrytning (vertikal sidbrytning) till vänster om den markerade cellen.  
En manuell kolumnbrytning känner du igen på den mörkblå vertikala linjen i tabellen.  
Infoga celler  
Här bestämmer du i en dialogruta vilka alternativ som ska gälla när nya celler infogas i dokumentet.  
Information om hur du kan radera celler får du på menyn Redigera - Radera celler.  
Urval  
I detta område kan Du välja på vilket sätt Du vill infoga celler i tabellen.  
Antal och position för de celler som ska infogas bestämmer Du genom att dessförinnan markera cellerna i tabellen.  
Flytta celler nedåt  
Med detta alternativ flyttas innehållet i cellerna i det markerade området nedåt när nya celler infogas.  
Flytta celler åt höger  
Med det här alternativet flyttar Du innehållet i cellerna i det markerade området åt höger när nya celler infogas.  
Infoga hela rader  
Markeringen i tabellen avgör infogningspositionen.  
Antalet rader som ska infogas bestäms av antalet markerade rader.  
Innehållen i de ursprungliga raderna förskjuts nedåt när nya rader infogas.  
Infoga hela kolumner  
Markeringen i tabellen avgör infogningspositionen.  
Antalet kolumner som ska infogas bestämms av antalet markerade kolumner.  
Innehållen i de ursprungliga kolumnerna förskjuts åt höger när nya kolumner infogas.  
Rader  
Med det här kommandot infogar du en ny rad i tabellen framför den aktiva cellen.  
Om flera rader är markerade när du väljer kommandot, infogas lika många rader som är markerade.  
De befintliga raderna förskjuts nedåt.  
Kolumner  
Med det här kommandot infogar du en ny kolumn i tabellen framför den aktiva kolumnen.  
Om flera kolumner är markerade när du väljer detta kommando infogas lika många kolumner som för tillfället är markerade.  
De befintliga kolumnerna förskjuts åt höger.  
Infoga tabell  
Här definierar du alternativen för att infoga en ny tabell.  
Du kan skapa en helt ny tabell eller skapa tabellen utifrån en fil, för att sedan infoga den i det aktuella tabelldokumentet.  
Position  
I detta område definierar du var tabellen ska infogas i dokumentet.  
Före aktuell tabell  
Med detta alternativ infogar du en ny tabell omedelbart före den aktuella tabellen.  
Efter aktuell tabell  
Med detta alternativ infogar du en ny tabell omedelbart efter den aktuella tabellen.  
Tabell  
I det här området definierar du om nya eller befintliga tabeller ska infogas i dokumentet.  
Skapa ny  
Med det här alternativet skapar du en ny tabell, som du kan ge ett namn i fältet Namn.  
Antal  
I detta rotationsfält kan du definiera antalet tabeller som ska infogas.  
Namn  
Här skriver du tabellens namn.  
Tabellnamn kan bestå av bokstäver och siffror.  
Skapa från fil  
Om du vill infoga ytterligare en tabell från en befintlig fil i det aktuella tabelldokumentet klickar du på det här alternativfältet.  
Genomsök  
Med den här kommandoknappen öppnar Du en dialogruta där Du kan välja en fil.  
Dialogrutan Infoga är i allt väsentligt densamma som dialogrutan Öppna på Arkiv -menyn.  
Valda tabeller  
Om Du har valt en fil med hjälp av knappen Genomsök visas den valda filens tabeller i listrutan.  
Under fältet visas filens sökväg.  
Markera den tabell som ska infogas i dokumentet i den här listrutan.  
Länka  
Om Du vill länka samman det aktuella dokumentet med den tabell som markerats i listrutan klickar Du här.  
Funktionsautopilot  
Här skapar du formler interaktivt med hjälp av Funktionsautopiloten.  
Innan du startar Funktionsautopiloten markerar du en cell eller ett cellområde där formeln ska infogas i den aktuella tabellen.  
Funktionsautopiloten innehåller två flikar:  
Under fliken Funktioner skapar du en formel, och under fliken Struktur granskar du formelns uppbyggnad.  
Fliken Funktioner  
Lista över kategorier och funktioner  
Kategori  
I det här kombinationsfältet ser du alla områden som funktionerna är indelade i.  
Om du väljer en kategori visas de tillhörande funktionerna i listrutan nedanför.  
Om du väljer "Senast använd" visas funktioner som redan har använts.  
Funktion  
I den här listrutan visas funktionerna i den valda kategorin.  
Välj en funktion genom att dubbelklicka på den.  
Om du klickar en gång visas en kort funktionsbeskrivning.  
Matris  
Om den här rutan är markerad, skapas en matris i det markerade tabellområdet, d.v.s. ett sammanhängande cellområde där den valda funktionen infogas som matrisformel.  
Varje cell i matrisen innehåller formeln, men inte som kopior utan som gemensam formel för alla celler i matrisen.  
Rutan Matris har samma funktion som tangentkombinationen Kommando Ctrl +Skift+Retur när du matar in och bekräftar en formel i tabellen: formeln infogas som matrisformel, vilket anges med två klammerparenteser.  
Den maximala storleken på ett matrisområde är 128 celler.  
Inmatningsområdet Argument  
När du väljer ut en funktion öppnas ett område på den högra sidan i Funktionsautopiloten där du kan ange argument.  
Om du ska välja en cellreferens som argument klickar du direkt på cellen, eller drar upp det önskade området i tabellen med nedtryckt musknapp.  
Numeriska och andra värden och referenser kan du också ange direkt i motsvarande fält i dialogrutan.  
Lägg märke till de särskilda regler som gäller när du anger datum.  
Klicka på OK så att resultatet förs in i tabellen.  
Delresultat  
När du anger argumenten i funktionen utförs beräkningen.  
I den här förhandsvisningen ser du om funktionsberäkningen kan utföras med de angivna argumenten.  
Om argumenten leder till ett fel, visas här motsvarande felkod.  
De inmatningar som är nödvändiga visas fetstilta med namn som står framför kommandoknappen.  
f( x) (beror av den valda funktionen)  
Genom att klicka på någon av de här kommandoknapparna går du en nivå djupare in i funktionsautopiloten.  
Du kan då använda den till att införa en funktion i stället för ett värde eller en referens i fältet bredvid kommandoknappen.  
Argument / Parameter / Cellreferens (beroende på vald funktion)  
Antalet textfält beror på funktionen.  
Du kan ange argument direkt i argumentfälten eller genom att klicka i en cell i tabellen.  
Resultat  
I det här förhandsvisningsfältet kan Du se resultatet av Dina beräkningar innan Du bekräftar dem med OK.  
Formel  
I det här fältet visas den skapade formeln.  
Här kan Du göra inmatningar direkt eller skapa formeln med hjälp av funktionsautopiloten.  
<<Tillbaka  
Med den här kommandoknappen går du till vänster i formelfönstret genom formelns beståndsdelar och markerar dem samtidigt.  
Om du vill markera en enskild funktion i en längre formel som består av flera funktioner, räcker det att dubbelklicka på funktionen i formelfönstret.  
Nästa >>  
Med den här kommandoknappen stegar Du åt höger genom formelkomponenterna i formelfönstret och ångrar därmed de markeringar som Du har gjort med kommandoknappen <<Tillbaka.  
Med knappen kan Du också föra över funktioner till formeln.  
Välj en funktion och klicka sedan på kommandoknappen.  
Den valda funktionen visas i formelfönstret.  
Om Du t ex vill ersätta de senaste två infogningarna med en ny funktion, klickar Du två gånger på kommandoknappen <<Tillbaka.  
Du kan ersätta det markerade formelområdet med en ny funktion genom att välja den och klicka på kommandoknappen Nästa>>.  
Du kan även föra över en funktion från urvalsfönstret genom att dubbelklicka.  
Avbryt  
Med den här kommandoknappen avslutar du funktionsautopiloten utan att överta någon formel.  
OK  
Med den här kommandoknappen avslutar du funktionsautopiloten och övertar formeln till den aktuella cellen eller cellerna.  
Lista över kategorier och funktioner  
Fliken Struktur  
Under den här fliken kan du se funktionsuppbyggnadens struktur.  
Om du startar Funktionsautopiloten medan cellmarkören står i en cell som redan innehåller en funktion, öppnas fliken Struktur där strukturen hos den aktuella formeln visas.  
Struktur  
Här visas funktionen hierarkiskt.  
Du kan öppna eller stänga formelposterna med plus - eller minustecknet när du vill se resp. dölja argumenten.  
De enskilda argumenten visas med en blå punkt om de är korrekt angivna.  
En röd punkt anger att datatypen är fel.  
Om Du t ex har angett en text som argument för funktionen SUMMA, visas argumentet i rött, eftersom den funktionen bara tillåter tal som argument.  
Kategorier och funktioner  
I det här avsnittet beskrivs funktionerna i %PRODUCTNAME Calc.  
De olika funktionerna är sammanfattade i praktiska kategorier i Funktionsautopiloten i %PRODUCTNAME Calc.  
Dessutom har du tillgång till operatorer.  
Databas  
Datum & Tid  
Finans  
Information  
Logisk  
Matematik  
Matris  
Statistik  
Tabell  
Text  
Add-In  
Här hittar Du de funktioner i %PRODUCTNAME Calc, som gäller hantering av data som sammanfattats radvis till dataposter.  
Funktionerna är följande:  
DANTAL, DANTALV, DHÄMTA, DMAX, DMIN, DMEDEL, DPRODUKT, DSTDAV, DSTDAVP, DSUMMA, DVARIANS, DVARIANSP.  
De beskrivs nedan.  
Öppna alltid sidan 2 i Funktionsautopiloten där Du kan jämföra den beskrivna funktionen.  
Kategorin Databas kan på grund av sitt namn förväxlas med en koppling till en databas i %PRODUCTNAME.  
Men det finns ingen som helst samband mellan en databas i %PRODUCTNAME och kategorin Databas i %PRODUCTNAME Calc.  
Titta på exempeltabellen som i området A1:E10 listar de barn som är inbjudna till Joes födelsedag.  
Därefter följer ålder (år), skolväg (m) och kroppsvikt (kg).  
A  
B  
C  
D  
E  
1  
Namn  
Klass  
Ålder  
Skolväg  
Vikt  
2  
Andy  
3  
9  
150  
40  
3  
Betty  
4  
10  
1000  
42  
4  
Charles  
3  
10  
300  
51  
5  
Daniel  
5  
11  
1200  
48  
6  
Eva  
2  
8  
650  
33  
7  
Frank  
2  
7  
300  
42  
8  
Greta  
1  
7  
200  
36  
9  
Hans  
3  
9  
1200  
44  
10  
Irene  
2  
8  
1000  
42  
11  
12  
13  
Namn  
Klass  
Ålder  
Skolväg  
Vikt  
14  
>600  
15  
16  
DANTAL  
5  
Formeln i cell B16 lyder =DANTAL( A1:E10;A1:E10;A13:E14)  
Parametrarna för samtliga databasfunktioner har följande betydelse:  
databas är det cellområde som definierar databasen.  
databasfält anger vilket databasfält som används för en relaterad referenshänvisning om en sådan är möjlig för databasfunktionen.  
Om Du vill referera till en kolumn genom namnet i kolumnhuvudet, sätter Du namnet inom citattecken.  
sökkriterier är det cellområde som innehåller sökkriterier.  
Om Du skriver flera kriterier på en rad, kopplas dessa kriterier ihop med OCH.  
Om Du skriver kriterier på olika rader under varandra, kopplas dessa kriterier ihop med ELLER.  
Tomma celler i sökkriteriernas område ignoreras.  
Under Verktyg - Alternativ - Tabelldokument - Beräkna kan du välja hur %PRODUCTNAME Calc ska hantera sökning efter exakta överensstämmelser.  
DANTAL  
DANTAL räknar antalet rader (dataposter) i en databas som överensstämmer med de inmatade sökkriterierna som innehåller numeriska värden.  
Syntax  
DANTAL( databas; databasfält; sökkriterier)  
Parametern får dock inte vara tom.  
Exempel  
I ovanstående exempel vill vi veta hur många barn som har en skolväg som överskrider 600 m.  
Resultatet ska sparas i cell B16.  
Placera markören i cell B16.  
Skriv formeln =DANTAL( A1:E10;A1:E10;A13:E14) i B16.  
Du kan även skriva formeln =DANTAL( A1:E10;0;A13:E14) (se syntax-anmärkning ovan).  
När Du anger områdena kan Du även ta hjälp av Funktionsautopiloten.  
databas är området med de data som ska utvärderas, inklusive deras huvuden, i det här fallet alltså A1:E10. databasfält definierar kolumnen för sökkriterierna, dvs skolväg (m) i detta fall. sökkriterier är det område där Du kan skriva in sökvillkoren.  
I det här fallet omfattar området A13:E14.  
Om Du t ex vill veta hur många barn i klass 2 som är äldre än 7 år, tar Du bort posten >600 i cell D14, anger sedan "2" i cell B14 under Klass och anger därefter ">7 "i cell C14.  
Resultatet är 2.  
Det finns två barn i klass 2 som är äldre än 7 år.  
Eftersom båda kriterierna står på samma rad, länkas de med ett logiskt OCH.  
ANTAL.TOMMA, ANTAL.OM.  
DANTALV  
DANTALV räknar antalet rader (dataposter) i en databas som överensstämmer med de inmatade sökkriterierna och som innehåller numeriska eller alfanumeriska värden.  
Syntax  
DANTALV( databas; databasfält; sökkriterier)  
Exempel  
I ovanstående exempel kan Du t ex söka efter det antal barn vars namn börjar på E eller någon därpå följande bokstav i alfabetet.  
Redigera formeln i B16 genom att komplettera funktionsnamnet DANTAL med bokstaven V.  
Ta bort de gamla sökkriterierna och ange "=E" under Namn i fält A14.  
Svaret är 5.  
Om Du nu t ex tar bort alla siffervärden för Greta, dvs på rad 8, ändras svaret till 4.  
Rad 8 räknas inte med längre eftersom den inte innehåller några värden (namnet Greta är bara text, inget värde).  
ANTAL.TOMMA, ANTAL.OM.  
DHÄMTA  
DHÄMTA fastställer innehållet i den ena cellen i en databas som det refereras till genom de inmatade sökkriterierna.  
Om det uppstår något fel returnerar funktionen #VÄRDE!, om ingen cell hittas, eller Err502 om flera celler hittas.  
Syntax  
DHÄMTA( databas; databasfält; sökkriterier)  
Exempel  
Vi vill i exemplet ovan ta reda på i vilken klass det barn går vars namn vi skriver in under Namn i cell A14.  
Dess lydelse skiljer sig något från de båda tidigare exemplen eftersom vi här bara får ange en kolumn (ett databasfält) för databasfält.  
Ange följande formel:  
=DHÄMTA( A1:E10; klass;A13:E14)  
Om Du nu skriver in namnet Frank i A14, får Du svaret 2.  
Frank går i 2:a klass.  
Du kan även skriva "ålder" i stället för "klass ", och får då Franks ålder.  
På rad 14 kan Du även välja att bara ange ett värde i cell C14, nämligen 11, och radera övriga poster på raden.  
Redigera formeln i B16 på följande sätt:  
=DHÄMTA( A1:E10 ;"namn";A13:E14)  
Nu frågar Du alltså efter namnet, och inte klassen.  
Svaret får Du direkt:  
Daniel är det enda barnet som är 11 år gammalt.  
DMAX  
DMAX fastställer det högsta värde som förekommer i en cell (datafält) på respektive rad (datapost) i en databas, och som överensstämmer med de inmatade sökkriterierna.  
Syntax  
DMAX( databas; databasfält; sökkriterier)  
Exempel  
Hur mycket väger det tyngsta barnet i varje klass?  
Ange följande formel i B16:  
=DMAX( A1:E10 ;"vikt";A13:E14)  
På rad 14 under Klass skriver Du nu i en följd 1, 2, 3 osv.  
Efter varje inmatning visas som resultat vikten för det tyngsta barnet i respektive klass.  
DMIN  
DMIN fastställer det lägsta värde som förekommer i en cell (datafält) på respektive rad (datapost) i en databas, och som överensstämmer med de inmatade sökkriterierna.  
Syntax  
DMIN( databas; databasfält; sökkriterier)  
Exempel  
Hur lång är den kortaste skolvägen för barnen i respektive klass?  
Ange följande formel i B16:  
=DMIN( A1:E10 ;"skolväg";A13:E14)  
På rad 14 under Klass skriver Du nu i en följd 1, 2, 3 osv.  
Efter varje inmatning visas som resultat skolvägens längd för det barn ur denna klass som har den kortaste skolvägen.  
DMEDEL  
DMEDEL fastställer medelvärdet för innehållet i alla celler (datafält) på alla rader (dataposter) i en databas som motsvarar de inmatade sökkriterierna.  
Syntax  
DMEDEL( databas; databasfält; sökkriterier)  
Exempel  
Hur stor är medelvikten för alla jämnåriga barn?  
Ange följande formel i B16:  
=DMEDEL( A1:E10 ;"vikt";A13:E14)  
På rad 14 under Ålder skriver Du nu i en följd 7, 8, 9 osv.  
Efter varje inmatning visas som resultat medelvikten för alla barn i den angivna åldern.  
DPRODUKT  
DPRODUKT multiplicerar ett databasfälts alla celler på alla rader (dataposter) i en databas som motsvarar de inmatade sökkriterierna.  
Syntax  
DPRODUKT( databas; databasfält; sökkriterier)  
Exempel  
När det gäller det ovanstående födelsedags-exemplet går det inte att använda den här funktionen på något meningsfullt sätt.  
DSTDAV  
Här behandlas dataposterna som ett stickprov.  
Vi vill alltså dra slutsatser utifrån "våra" barn för alla barn (vilket givetvis inte ger några tillförlitliga resultat om underlaget inte är mer än något tusentals barn).  
Syntax  
DSTDAV( databas; databasfält; sökkriterier)  
Exempel  
Hur hög är standardavvikelsen när det gäller vikten för barn i en viss ålder?  
Ange följande formel i B16:  
=DSTDAV( A1:E10 ;"vikt";A13:E14)  
På rad 14 under Ålder skriver Du nu i en följd 7, 8, 9 osv.  
Efter varje inmatning visas som resultat standardavvikelsen för vikten för alla barn i den angivna åldern.  
DSTDAVP  
DSTDAVP bestämmer standardavvikelsen för ett databasfälts alla celler på alla rader (dataposter) i en databas som motsvarar de inmatade sökkriterierna.  
Vi vill alltså bara dra slutsatser om våra barn, inte om andra barn för vilka vi inte har samlat in några data.  
Syntax  
DSTDAVP( databas; databasfält; sökkriterier)  
Exempel  
Hur hög är standardavvikelsen för vikten för alla jämnåriga barn på Joes födelsedagskalas?  
Ange följande formel i B16:  
=DSTDAVP( A1:E10 ;"vikt";A13:E14)  
På rad 14 under Ålder skriver Du nu i en följd 7, 8, 9 osv.  
Efter varje inmatning visas som resultat standardavvikelsen för vikten för alla barn i den angivna åldern som vi har vägt.  
DSUMMA  
DSUMMA bestämmer summan för ett databasfälts alla celler i en databas på alla rader (dataposter) som motsvarar de inmatade sökkriterierna.  
Syntax  
DSUMMA( databas; databasfält; sökkriterier)  
Exempel  
Hur lång är den totala skolvägen för alla barn på Joes födelsedagskalas som går i 2:a klass?  
Ange följande formel i B16:  
=DSUMMA( A1:E10 ;"skolväg";A13:E14)  
På rad 14 under Klass skriver Du nu enbart 2.  
Som resultat visas summan av skolvägarna för alla barn ur 2:a klass, nämligen 1950.  
SUMMA.OM  
DVARIANS  
Här behandlas dataposterna som ett stickprov.  
Vi vill alltså dra slutsatser utifrån "våra" barn för alla barn (vilket givetvis inte ger några tillförlitliga resultat om underlaget inte är mer än något tusentals barn).  
Syntax  
DVARIANS( databas; databasfält; sökkriterier)  
Exempel  
Hur hög är variansen för vikten för alla jämnåriga barn?  
Ange i B16 denna formel:  
=DVARIANS( A1:E10 ;"vikt";A13:E14)  
På rad 14 under Ålder skriver Du nu i en följd 7, 8, 9 osv.  
Efter varje inmatning visas som resultat variansen för vikten för alla barn i den angivna åldern.  
DVARIANSP  
DVARIANSP bestämmer variansen för ett databasfälts alla celler i en databas på alla rader (dataposter) som motsvarar de inmatade sökkriterierna.  
Vi vill alltså bara dra slutsatser om våra barn, inte om andra barn för vilka vi inte har samlat in några data.  
Syntax  
DVARIANSP( databas; databasfält; sökkriterier)  
Exempel  
Hur hög är variansen för vikten för alla jämnåriga barn på Joes födelsedagskalas?  
Ange följande formel i B16:  
=DVARIANSP( A1:E10 ;"vikt";A13:E14)  
På rad 14 under Ålder skriver Du nu i en följd 7, 8, 9 osv.  
Efter varje inmatning visas som resultat variansen för vikterna för alla barn i den angivna åldern på Joes födelsedagskalas.  
Kategori Datum & Tid  
Här hittar du de %PRODUCTNAME Calc-funktioner som infogar och redigerar datum och klockslag.  
Det rör sig om funktionerna ARBETSDAGAR, DAG, DAGAR, DAGAR360, DATUM, DATUMVÄRDE, EDATUM, IDAG, KLOCKSLAG, MINUT, MÅNAD, NETTOARBETSDAGAR, NU, PÅSKDAGEN, SEKUND, SLUTMÅNAD, TIDVÄRDE, TIMME, VECKODAG, VECKONR, VECKONR_ADD, ÅR och ÅRDEL.  
De beskrivs nedan.  
Du kan jämföra den beskrivna funktionen genom att öppna sidan 2 i Funktionsautopiloten.  
%PRODUCTNAME behandlar internt datum - / tidsvärden som numeriska värden.  
12:00 om till 36526,50.  
Värdet framför kommat motsvarar datumet och värdet efter kommat tiden.  
Om du skulle råka konfronteras med sådana numeriska framställningar av datum och tid bör du kontrollera att rätt talformat (datum eller tid) har ställts in.  
Markera den cell som innehåller datum - / tidsvärdet och välj Formatera celler... på snabbmenyn.  
Under fliken Tal hittar du funktionerna för att bestämma talformatet.  
Under Verktyg - Alternativ - %PRODUCTNAME - Allmänt finns området Tvåsiffriga årtal.  
Där ställer du in tidsperioden då tvåsiffriga årtal ska gälla.  
Observera att ändringar som du gör här påverkar en del av följande funktioner.  
Observera följande när du arbetar med datumangivelser: om du använder bindestreck och snedstreck som skiljetecken i en formel tolkas det som del av en formel och inte som datum.  
Om du anger 20 / 07 / 54 eller 54-07-20 i stället för 54.07.20 leder det till ett felaktigt resultat.  
Sätt därför datum med snedstreck eller bindestreck inom citattecken, t.ex. "54-07-20".  
ARBETSDAGAR  
Resultatet är ett datumtal som kan formateras som datum.  
Du ser då datumet på en dag som ligger ett visst antal Arbetsdagar före eller efter ett Startdatum.  
Syntax  
ARBETSDAGAR( Startdatum;Dagar;Lediga dagar)  
Startdatum: datumet från vilket beräkningen sker.  
Om startdatumet är en arbetsdag räknas den dagen med.  
Dagar: antalet arbetsdagar.  
Positivt värde för ett resultat efter startdatum, negativt värde för ett resultat före startdatum.  
Lediga dagar: valfri lista med lediga dagar.  
Det är dagar då man inte arbetar.  
Ange ett cellområde där de lediga dagarna är listade en och en.  
Exempel  
Vilket datum är det 17 arbetsdagar efter den 1 december 2001?  
Startdatumet "2001-12-01" står i C3, antalet arbetsdagar står i D3.  
I cellerna F3 till J3 står följande lediga dagar vid jul och nyår: "2001-12-24", "2001-12-25", "2001-12-26", "2001-12-31", "2002-01-01".  
=ARBETSDAGAR( C3;D3;F3:J3) ger resultatet 01-12-28.  
Formatera det seriella datumtalet som datum.  
ÅRDEL  
Resultatet är ett tal mellan 0 och 1 som representerar bråkdelen av ett år mellan Startdatum och Slutdatum.  
Syntax  
ÅRDEL( Startdatum;Slutdatum;Bas)  
Startdatum och slutdatum: två datumvärden.  
Bas: valfritt, anger hur året ska beräknas.  
Bas  
Beräkning  
0 eller saknas  
US-metod (NASD), 12 månader om 30 dagar  
1  
exakt antal dagar per månad, exakt antal dagar per år  
2  
exakt antal dagar per månad, år har 360 dagar  
3  
exakt antal dagar per månad, år har 365 dagar  
4  
Europa-metod, 12 månader om 30 dagar  
Exempel  
Vilken bråkdel av året 2001 ligger mellan 2002-01-01 och 2001-07-01?  
=ÅRDEL( "2002-01-01"; "2002-07-01";1) ger resultatet 0,495890.  
DATUM  
Den här funktionen omvandlar ett datum, skrivet som år, månad, dag, till ett internt tal och visar det i cellens formatering.  
Då visas datumets interna tal som ett tal.  
Syntax  
DATUM( år; månad; dag)  
år är ett heltal mellan 1583 och 9956 eller 0 och 29.  
Under Verktyg - Alternativ - %PRODUCTNAME - Allmänt kan du ställa in från vilket årtal ett tvåsiffrigt tal ska identifieras som 20xx.  
månad är ett tal mellan 1 och 12 med vilket månadstalet anges.  
dag är ett tal mellan 1 och 31, som fastställer dagen i månaden.  
Om värdena för månad och dag är större avräknas de med spill till nästa decimal.  
Om Du skriver =DATUM( 00;12;31), får Du som resultat 2000-12-31.  
Om Du skriver =DATUM( 00;13;31) får Du det korrekta 2001-01-31.  
Som argument i funktionen DATUM kan Du skriva in datumuppgifter direkt eller göra områdesreferenser.  
Exempel  
DATUM( "00;1;1") ger 2000-01-01  
DATUMVÄRDE, IDAG, ÅR, NU, MÅNAD, DAG, TIDVÄRDE.  
DATUMVÄRDE  
DATUMVÄRDE beräknar det interna datumtalet ur en text som Du anger inom citattecken och som representerar ett möjligt inmatningsformat för datum.  
Det interna talet, som anges som ett naturligt tal, får Du ur det datumsystem som används i %PRODUCTNAME för beräkning av datumuppgifter.  
Syntax  
DATUMVÄRDE( "text")  
text är ett giltigt datumuttryck som måste anges inom citattecken.  
Exempel  
DATUMVÄRDE( "54.7.20") ger 19925  
IDAG, NU, TIDVÄRDE.  
EDATUM  
Resultatet är ett datum som ligger ett antal Månader före eller efter Startdatum.  
Det är bara månader som räknas, inte dagar.  
Syntax  
EDATUM( Startdatum;Månader)  
Startdatum: ett datum.  
Månader: antalet månader.  
Exempel  
Vilket datum är det en månad före 2001-03-31?  
=EDATUM( "2001-03-31";-1) ger resultatet 2001-02-28.  
IDAG  
Infogar det aktuella datumet i datorn.  
Värdet uppdateras när Du öppnar dokumentet igen, eller när dokumentets värdeintervall ändras.  
Syntax  
IDAG()  
Idag är en funktion utan argument.  
Exempel  
IDAG() ger det aktuella datumet i datorns systemklocka i formen 2000-02-02.  
DATUM, NU, DAG.  
ÅR  
Beräknar för ett tal det år som tilldelats enligt den interna uträkningen.  
Syntax  
ÅR( tal)  
tal anger det interna datumvärde för vilket årtalet ska beräknas.  
Exempel  
ÅR( 1) ger 1899  
ÅR( 2) ger 1900  
ÅR( 33333,33) ger 1991  
IDAG, NU, MINUT, MÅNAD, SEKUND, TIMME, DAG, VECKODAG.  
NU  
Anger datum och klockslag i enlighet med datorns systemklocka.  
Värdet uppdateras om Du beräknar dokumentet på nytt eller varje gång som cellvärdet ändras.  
Syntax  
NU()  
Exempel  
=NU( )-A1 ger differensen mellan datumet i A1 och nu.  
Formatera resultatet som tal.  
DATUM, ÅR, MINUT, MÅNAD, TIMME, DAG, VECKODAG.  
VECKONR  
VECKONR beräknar årets kalendervecka för det interna datumvärdet.  
Syntax  
VECKONR( tal; läge)  
tal är det interna datumtalet.  
läge beräknar när veckan börjar och typ av beräkning.  
1 = Söndag  
2 = Måndag  
Exempel  
VECKONR( "95.1.1";1) returnerar 1 (den 1 / 1 95 var en söndag)  
VECKONR( "95.1.1";2) returnerar 52 (om veckan börjar med måndag hör denna söndag till sista veckan på det föregående året).  
VECKONR_ADD  
Resultatet är numret på kalenderveckan till ett Datum.  
Syntax  
VECKONR_ADD( Datum;Returtyp)  
Datum: datumet inom kalenderveckan.  
Returtyp:  
1 om veckan början på söndagar, 2 om veckan börjar på måndagar.  
Exempel  
I vilken kalendervecka ligger 2001-12-24?  
=VECKONR_ADD( "2001-12-24";1) ger resultatet 52.  
MINUT  
MINUT beräknar antalet minuter till det interna tidvärdet.  
Minutvärdet anges som ett tal mellan 0 och 59.  
Syntax  
MINUT( tal)  
tal är som tidvärde ett decimaltal för vilket antal minuter ska beräknas.  
Exempel  
MINUT( 8,999) returnerar 58  
MINUT( 8,9999) returnerar 59  
MINUT( NU()) returnerar det aktuella antalet minuter.  
ÅR, NU, MÅNAD, SEKUND, TIMME, DAG, VECKODAG.  
MÅNAD  
Beräknar månaden för det givna datumvärdet.  
Månaden anges som ett tal mellan 1 och 12.  
Syntax  
MÅNAD( tal)  
tal är som tidvärde ett decimaltal för vilket månaden ska beräknas.  
Exempel  
MÅNAD( NU)()) ger aktuell månad  
MÅNAD( C4) ger 7, när innehållet i C4 = 2000-07-07.  
ÅR, NU, MINUT, TIMME, DAG, VECKODAG.  
SLUTMÅNAD  
Resultatet är datumet på den sista dagen i en månad som ligger ett visst antal Månader före eller efter Startdatum.  
Syntax  
SLUTMÅNAD( Startdatum; Månader)  
Startdatum: från detta datum sker beräkningen.  
Månader: månaden ska ligga så många månader före (negativt) eller senare (positivt).  
Exempel  
Vilken är den sista dagen i månaden som ligger 6 månader före den 12 september 2001?  
=SLUTMÅNAD( "2001-09-12";6) ger resultatet 2002-03-31.  
NETTOARBETSDAGAR  
Resultatet är antalet arbetsdagar mellan Startdatum och Slutdatum.  
Lediga dagar kan dras ifrån.  
Syntax  
NETTOARBETSDAGAR( Startdatum;Slutdatum;Lediga dagar)  
Startdatum: datumet från vilket beräkningen sker.  
Om startdatum är en arbetsdag räknas den dagen med.  
Slutdatum: datumet fram till vilket beräkningen sker.  
Om slutdatum är en arbetsdag räknas den dagen med.  
Det är dagar när man inte arbetar.  
Ange ett cellområde där de lediga dagarna är listade en och en.  
Exempel  
Hur många arbetsdagar är det mellan 2001-12-15 och 2002-01-15?  
Startdatumet står i C3, slutdatumet står i D3.  
I cellerna F3 till J3 står följande lediga dagar till jul och nyår: "2001-12-24", "2001-12-25", "2001-12-26", "2001-12-31", "2002-01-01".  
=NETTOARBETSDAGAR( C3;D3;F3:J3) ger resultatet 17 arbetsdagar.  
PÅSKDAGEN  
Beräknar för ett visst givet år det datum som påsksöndagen infaller på.  
År är ett heltal från 1583 till 9956 (ifall ingen kalenderreform kommer innan dess), respektive 0 till 99.  
Funktionen ger det interna datumtalet för påskdagen det aktuella året Påskdagen är den första söndagen efter den första fullmånen efter vårdagjämningen.  
Du kan beräkna ytterligare rörliga helgdagar genom att göra en enkel addition med detta datum:  
Annandag påsk = PÅSKDAGEN() + 1  
Långfredagen = PÅSKDAGEN() - 2  
Pingstdagen = PÅSKDAGEN() + 49  
Annandag pingst = PÅSKDAGEN() +50  
Exempel  
PÅSKDAGEN( 2000) ger den 2000-04-23  
PÅSKDAGEN( 2000 )+49 returnerar det interna värdet 36688.  
Om du formaterar det med datumformatet TTMMJJJJ får du 2000-06-11.  
SEKUND  
Beräknar sekunden för det givna tidvärdet.  
Sekundvärdet anges som ett tal mellan 0 och 59.  
Syntax  
SEKUND( tal)  
tal är som tidvärde ett decimaltal för vilket sekunden ska beräknas.  
Exempel  
SEKUND( NU()) ger aktuell sekund  
SEKUND( C4) ger 17, när innehållet i C4 = 12:20:17.  
DATUM, ÅR, NU, MINUT, MÅNAD, TIMME, DAG, VECKODAG.  
TIMME  
Beräknar timmen till det givna tidvärdet.  
Timmen anges som ett tal mellan 0 och 23.  
Syntax  
TIMME( tal)  
tal är som tidvärde ett decimaltal för vilket timmen ska beräknas.  
Exempel  
TIMME( NU()) ger aktuell timme  
TIMME( C4) ger 17, när innehållet i C4 = 17:20:00.  
ÅR, NU, MINUT, MÅNAD, DAG, VECKODAG.  
DAG  
Beräknar dagen för det givna datumvärdet.  
Dagen anges som ett tal mellan 1 och 31.  
Du kan också använda negativt datum / negativ tid för beräkningar.  
Syntax  
DAG( tal)  
tal är som tidvärde ett decimaltal för vilket dagen ska beräknas.  
Exempel  
DAG( 1) ger 31 (eftersom %PRODUCTNAME börjar räkna vid noll den 31 / 12 1899)  
DAG( NU()) ger dagen idag.  
DAG( C4) ger 5, när innehållet i C4 = 1901-08-05.  
IDAG, ÅR, NU, MINUT, MÅNAD, SEKUND, TIMME, VECKODAG.  
DAGAR  
Beräknar differensen mellan två datumtal.  
Resultatet är ett heltal och anger antal dagar mellan de två datumen.  
Syntax  
DAGAR( datum_2;datum_1)  
datum_1 är det senare datumet, datum_2 är det tidigare datumet.  
Om Du anger datumtalen i omvänd ordningsföljd får funktionen ett negativt tal som resultat.  
Exempel  
DAGAR( "2010.1.1"; NU()) ger antalet dagar från idag och till den 1 januari 2010.  
DAGAR( "1990.10.10"; "1980.10.10") ger 3652.  
DAGAR360  
Beräknar differensen mellan två datumtal på basen 360 dagar per år, vilket är vanlig vid ränteberäkningar.  
Resultatet anges i form av ett heltal.  
Syntax  
DAGAR360( datum_1;datum_2;typ)  
Om datum2 ligger före datum1 i tiden får funktionen ett negativt tal som resultat.  
Den valfria parametern typ bestämmer typen av differensbildning.  
Om typ = 0 eller om parametern saknas används den amerikanska metoden (NASD, National Association of Securities Dealers).  
Om typ <> 0 används den europeiska metoden.  
Här får Du ytterligare information om DAGAR360.  
Exempel  
DAGAR360( 00.01.01; NU()) ger antalet räntedagar från den 1:e detta år och fram till idag.  
DAG.  
VECKODAG  
Beräknar veckodagen för det givna datumvärdet.  
Veckodagen anges som ett tal mellan 1 och 7 (vid typ=3 som ett tal mellan 0 och 6).  
1 är lika med söndag, såvida Du inte anger någon annan typ eller typ=1.  
När typ=2 börjar räkningen med måndag=1, när typ=3 börjar räkningen med måndag=0.  
Syntax  
VECKODAG( tal;typ)  
tal är som datumvärde ett decimaltal för vilket veckodagen ska beräknas.  
typ bestämmer typen av beräkning.  
För typ=1 gäller att veckodagarna räknas från och med söndag (detta är förinställt, även om parametern typ saknas), för typ=2 gäller att veckodagarna räknas från och med måndag=1, för typ=3 räknas veckodagarna från måndag=0.  
Dessa värden gäller bara för standarddatumformatet som du kan välja under Verktyg - Alternativ - Tabelldokument - Beräkna.  
Exempel  
VECKODAG( "2000.6.14") ger 4 (parametern typ saknas, därför gäller standardräkningen.  
Vid standardräkningen är söndag dagen med nummer 1.  
Den 14 / 6 2000 var en onsdag, alltså den fjärde dagen i veckan).  
VECKODAG( "1996.7.24"; 2) ger 3 (parametern typ är 2, alltså gäller att måndag är dagen med nummer 1.  
Den 24 / 7 96 är en onsdag, den har därför nummer 3).  
VECKODAG( "24.7.1996"; 1) ger 4 (parametern typ är 1, alltså gäller att söndag är dagen med nummer 1.  
Den 24 / 7 1996 är en onsdag, den har därför nummer 4).  
VECKODAG( NU()) ger numret för dagens veckodag.  
Om du vill veta om en dag som står i A1 är en arbetsdag eller inte, använder du funktionerna OM och VECKODAG så här:  
OM( VECKODAG(A1;2)<6 ;"Arbetsdag" ;"Veckoslut")  
IDAG, NU, DAG, TEXT.  
KLOCKSLAG  
KLOCKSLAG beräknar det aktuella tidvärdet ur värden för timmar, minuter och sekunder.  
Du kan använda funktionen för att ur dessa tre enskilda beståndsdelar räkna om en tidsangivelse till ett decimalt tidvärde.  
Syntax  
KLOCKSLAG( timme; minut; sekund)  
Timme förinmatas med ett heltal.  
Minut förinmatas med ett heltal.  
Sekund förinmatas med ett heltal.  
Exempel  
KLOCKSLAG( "0;0;0") ger 00:00:00  
KLOCKSLAG( "4;20;4") ger 04:20:04  
NU, MINUT, SEKUND, TIMME.  
TIDVÄRDE  
TIDVÄRDE beräknar det interna tidtalet ur en text som anges inom citattecken och som representerar ett möjligt inmatningsformat för tid.  
Det interna talet, som anges som ett decimaltal, är ett resultat av det datumsystem som används i %PRODUCTNAME för beräkning av datumuppgifter.  
Syntax  
TIDVÄRDE( "text")  
text är ett giltigt tidsuttryck som ska anges inom citattecken.  
Exempel  
Om du formaterar i tidsformatet HH:MM:SS får du 16:00:00.  
Om du formaterar med tidsformatet TT:MM:SS får du midnatt, d.v.s.  
DATUMVÄRDE, NU, MINUT, SEKUND, TIMME, KLOCKSLAG.  
Kategori Finans del 1  
I den här kategorin finns de finansmatematiska funktionerna i %PRODUCTNAME Calc.  
Funktionerna är följande:  
AMORDEGRC, AMORLINC, BELOPP, DB, DEGAVSKR, DISK, EFFRÄNTA, EFFRÄNTA_ADD, IR, LÖPTID_ADD, NUVÄRDE, RALÅN, UPPLOBLRÄNTA, UPPLRÄNTA och ÅRSAVSKR.  
Till finansfunktionerna del 2  
Till finansfunktionerna del 3  
AMORDEGRC  
Beräknar avskrivningsbeloppet för en avräkningsperiod som degressiv amortering.  
I motsats till AMORLINC används här en avskrivningskoefficient som beror på tillgångarnas livslängd.  
Syntax  
AMORDEGRC( Kostnader;Datum;Första period;Restvärde;Period;Ränta;Bas)  
Kostnader: anskaffningskostnaderna.  
Datum: anskaffningsdatumet.  
Första period: datumet för slutet på den första perioden.  
Restvärde: restvärde för tillgången i slutet av livslängden.  
Period: avräkningsperioden.  
Ränta: avskrivningssatsen.  
AMORLINC  
Beräknar avskrivningsbeloppet för en avräkningsperiod som linjär amortering.  
Om tillgången köps in under avräkningsperioden tas det proportionella avskrivningsbeloppet med i beräkningen.  
Syntax  
AMORLINC( Kostnader;Datum;Första period;Restvärde;Period;Ränta;Bas)  
Kostnader: anskaffningskostnader.  
Datum: anskaffningsdatum.  
Första period: datumet för slutet på den första avräkningsperioden.  
Restvärde: restvärdet för tillgången i slutet av livslängden.  
Period: avräkningsperioden.  
Ränta: avskrivningssatsen.  
UPPLRÄNTA  
Beräknar de upplupna räntorna för ett värdepapper med periodiska betalningar.  
Syntax  
UPPLRÄNTA( Emission;Första kupongdatum;Betalning;Nominell ränta;Nominellt värde;Frekvens;Bas)  
Emission: värdepapperets utgivningsdatum.  
Första kupongdatum: värdepapperets första räntedatum.  
Betalning: datumet för vilket de hittills upplupna räntorna ska beräknas.  
Nominell ränta: den årliga nominella räntan (kupongränta).  
Nominellt värde: värdepapperets nominella värde.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper ges ut den 28 februari 2001.  
Det första räntedatumet är den 31 augusti 2001.  
Betalningsdatumet är den 1 maj 2001.  
Nominell ränta är 0,1 eller 10%, det nominella värdet 1000 valutaenheter.  
Räntorna betalas halvårsvis (frekvens är 2).  
Bas är US-metoden (0) Hur höga är de upplupna räntorna?  
=UPPLRÄNTA( "2001-02-28"; "2001-08-31"; "2001-05-01"; 0,1; 1000; 2; 0) ger resultatet 16,94444.  
UPPLOBLRÄNTA  
Beräknar ett värdepappers upplupna räntor som betalas ut på förfallodagen.  
Syntax  
UPPLOBLRÄNTA( Emission;Betalning;Nominell ränta;Nominellt värde;Bas)  
Emission: värdepapperets utgivningsdatum.  
Betalning: förfallodagen.  
Nominell ränta: den årliga nominella räntan (kupongränta).  
Nominellt värde: värdepapperets nominella värde.  
Exempel  
Ett värdepapper ges ut den 1 april 2001.  
Förfallodagen är den 15 juni 2001.  
Nominell ränta är 0,1 eller 10%, det nominella värdet är 1000 valutaenheter.  
Hur höga är de upplupna räntorna?  
=UPPLOBLRÄNTA( "2001-04-01"; "2001-06-15"; 0,1; 1000; 3) ger resultatet 20,54795.  
BELOPP  
Beräknar beloppet som betalas ut vid en viss tidpunkt för ett värdepapper med fast ränta.  
Syntax  
BELOPP( Betalning;Förfallodag;Investering;Diskonteringsränta;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Investering: det investerade beloppet.  
Diskonteringsränta: den procentuella diskonteringen vid köpet av värdepapperet.  
Exempel  
Betalning:  
15 februari 1999, Förfallodag:  
15 maj 1999, Investering:  
1000 valutaenheter, Diskonteringsränta:  
5,75 procent, Bas: faktisk / 360 = 2.  
Beloppet som betalas ut på förfallodagen beräknas på följande sätt:  
=BELOPP( "1999-02-15" ;"1999-05-15";1000; 0,0575;2) returnerar 1014,420266.  
NUVÄRDE  
Beräknar det nuvarande värdet av en följd av regelbundna betalningar.  
Du kan använda den här funktionen till att beräkna hur stort belopp Du måste investera i dag för att det ska räcka till utbetalning av ett visst belopp (annuitet) vid ett visst antal utbetalningar.  
Du kan om Du vill ange hur mycket pengar som ska återstå när alla utbetalningar har gjorts.  
Du kan även ange om utbetalningen ska göras i början eller slutet av varje period.  
Du anger värdena som tal, uttryck eller referenser.  
Om Du t ex erhåller 8% i ränta varje år men skulle vilja ange månad som period, skriver Du 8% / 12 i fältet ränta. %PRODUCTNAME Calc beräknar automatiskt den korrekta faktorn.  
Syntax  
NUVÄRDE( ränta; Perioder; Betalning; Slutvärde; F)  
Ränta är räntesatsen för en periods betalning.  
Perioder är betalningstiden angiven i antalet perioder.  
Betalning är betalningen för en period.  
Slutvärde (valfritt) är det framtida värdet som ska bli över när alla betalningar är gjorda.  
F (valfritt) är förfallotidpunkten.  
F = 1 om betalningen görs under periodens början; F = 0 (standardvärde) om den görs vid dess slut.  
Exempel  
Hur högt är nuvärdet av en investering om 500 valutaenheter betalas ut varje månad och räntesatsen är 8% per år?  
Betalningstiden är 48 månader och som slutvärde ska 20 000 valutaenheter återstå.  
NUVÄRDE( 8% / 12;48;500;20000) = -35 019,37 valutaenheter.  
Med de givna förutsättningarna måste du alltså i dag betala 35 019,37 valutaenheter, om du vill erhålla 500 valutaenheter under 48 månader och vid periodens slut fortfarande ha 20 000 valutaenheter kvar.  
En moträkning visar att du kommer att få ut 48*500 valutaenheter + 20 000 valutaenheter = 44 000 valutaenheter.  
Skillnaden jämfört med det inbetalda beloppet 35 000 valutaenheter utgörs av de räntor som du kan tillgodoräkna dig.  
Tänk på att referenserna till konstanter ska vara absoluta referenser.  
Avskrivningsfunktionerna är ett exempel på den här typen av användning.  
AMORT, BETALNING, RÄNTA, RBETALNING, SLUTVÄRDE, PERIODER.  
ÅRSAVSKR  
Beräknar den digitala (aritmetiskt degressiva) avskrivningen.  
Den här funktionen använder Du för att beräkna avskrivningsdelen för en period i den totala avskrivningstiden för ett objekt.  
Vid digital avskrivning minskas avskrivningssumman från period till period med ett konstant belopp.  
Syntax  
ÅRSAVSKR( AV;RV;LL;TP)  
AV är tillgångens anskaffningsvärde.  
RV är tillgångens restvärde vid livslängdens slut.  
LL är livslängden uttryckt i antalet avskrivningsperioder.  
TP är den tidsperiod för vilken avskrivningen ska beräknas.  
Exempel  
En videoanläggning med ett anskaffningsvärde på 50 000 valutaenheter ska skrivas av årligen under fem år.  
Restvärdet ska vara 10 000 valutaenheter.  
Avskrivningen ska beräknas för det första året.  
ÅRSAVSKR( 50000;10000;5;1) = 13 333,33 valutaenheter.  
Avskrivningsbeloppet det första året är 13 333,33 valutaenheter.  
Du bör helst skapa en avskrivningstabell, så att Du lätt kan se avskrivningarna per tidsperiod.  
Om Du skriver in de olika avskrivningsformlerna i %PRODUCTNAME Calc ser Du också vilken form av avskrivning som är den lämpligaste i det här fallet.  
Fyll i tabellen enligt nedan:  
A  
B  
C  
D  
E  
1  
Anskaffningsvärde  
Restvärde  
Livslängd  
Tidsperiod  
ÅRSAVSKR  
2  
50 000 valutaenheter  
10 000 valutaenheter  
5  
1  
13 333,33 valutaenheter  
3  
2  
10 666,67 valutaenheter  
4  
3  
8 000,00 valutaenheter  
5  
4  
5 333,33 valutaenheter  
6  
5  
2 666,67 valutaenheter  
7  
6  
0,00 valutaenheter  
8  
7  
-  
9  
8  
-  
10  
9  
-  
11  
10  
-  
12  
13  
>0  
Summa  
40 000,00 valutaenheter  
Formeln i E2 lyder som följer:  
=ÅRSAVSKR( $A$2;$B$2;$C$2;D2)  
Den här formeln dupliceras i kolumn E till E10 (markera E2 och dra sedan nedåt i det nedre högra hörnet med musen).  
I cell E13 står den formel som kontrollsummerar alla avskrivningsbelopp.  
Du använder funktionen SUMMA.OM, eftersom de negativa värdena i E8:E11 inte får påverka resultatet.  
Villkoret >0 står i cell A13.  
Formeln i E13 lyder som följer:  
=SUMMA.OM( E2:E11;A13)  
Nu kan du se hur det blir om avskrivningstiden är 10 år, eller om restvärdet ska vara 1 valutaenhet, eller också anger du ett annat anskaffningsvärde och så vidare.  
DEGAVSKR, LINAVSKR, VDEGRAVSKR.  
DISK  
Beräknar diskonteringsräntan för ett värdepapper i procent.  
Syntax  
DISK( Betalning;Förfallodag;Pris;Inlösningsvärde;Bas)  
Betalning: datumet för värdepappersköpet.  
Förfallodag: datumet då värdepapperet förfaller.  
Pris: värdepapperets pris per 100 valutaenheter nominellt värde.  
Inlösningsvärde: värdepapperets inlösningsvärde per 100 valutaenheter nominellt värde.  
Exempel  
Ett värdepapper köps den 25 januari 2001; förfallodagen är den 15 november 2001.  
Hur hög är diskonteringsräntan vid faktisk / 365 beräkning (bas 3)?  
=DISK( "2001-01-25"; "2001-11-15"; 97; 100; 3) returnerar 0,03840 eller 3,84 procent.  
LÖPTID_ADD  
Beräknar löptiden för ett värdepapper med periodisk räntebetalning.  
Syntax  
LÖPTID_ADD( Betalning;Förfallodag;Nominell ränta;Avkastning;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Nominell ränta: den årliga nominella räntan (kupongränta).  
Avkastning: den årliga avkastningen för värdepapperet.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 1 januari 2001; förfallodagen är den 1 januari 2006.  
Avkastningen uppgår till 9,0%.  
Hur lång är löptiden vid faktisk / 365 beräkning (bas 3)?  
=LÖPTID_ADD( "2001-01-01"; "2006-01-01"; 0,08; 0,09; 2; 3)  
EFFRÄNTA  
Beräknar den årliga effektiva räntan utgående från en normalränta.  
I praktiken betalas normalräntan alltså i praktiken i förväg, och därigenom ökas den effektiva räntan med räntebetalningarna.  
Syntax  
EFFRÄNTA( NR;P)  
NR är nominalräntan.  
P är antalet periodiska räntebetalningar per år.  
Exempel  
Om nominalräntan per år är 9,75% och räntan ska betalas fyra gånger, hur hög blir då den verkliga räntan (effektivräntan)?  
Den årliga effektiva räntan är alltså 10,11%.  
NOMRÄNTA.  
EFFRÄNTA_ADD  
Beräknar den årliga effektiva räntan baserat på den nominella räntan och antalet räntebetalningar per år.  
Syntax  
EFFRÄNTA_ADD( Nominell ränta;Perioder)  
Nominell ränta: den årliga nominella räntan.  
Perioder: antalet räntebetalningar per år.  
Exempel  
Vad uppgår den effektiva räntan till vid 5,25% nominell ränta och kvartalsvis betalning?  
=EFFRÄNTA_ADD( 0,0525; 4) returnerar 0,053543 eller 5,3534%.  
DEGAVSKR  
Beräknar avskrivningen enligt den aritmetisk-degressiva metoden för en viss avskrivningsperiod.  
Den här avskrivningsformen använder Du när Du vill att avskrivningsvärdet ska vara störst i början av avskrivningen (i motsats till linjär avskrivning).  
Avskrivningsvärdet minskar för varje avskrivningsperiod med de avskrivningar som redan har dragits av från anskaffningsvärdet.  
Exempel är personbilar och IT-utrustning.  
Lägg märke till att bokföringsvärdet med den här beräkningsformen aldrig kan gå ner till noll.  
Syntax  
DEGAVSKR( AV;RV;LL;P;FA)  
AV är tillgångens anskaffningsvärde.  
RV är tillgångens restvärde vid livslängdens slut.  
LL är livslängden uttryckt i antalet avskrivningsperioder.  
P är periodlängden.  
FA (valfritt) är avskrivningsfaktorn.  
Om inget annat anges används faktorn 2.  
Exempel  
Ett datorsystem med ett anskaffningsvärde på 75 000 valutaenheter ska skrivas av månatligen under fem år.  
Restvärdet ska vara 1 valutaenhet.  
Faktorn är 2.  
DEGAVSKR( 75000;1;60;12;2) = 1 721,81 valutaenheter.  
Följaktligen är den degressiva avskrivningen den första månaden efter anskaffningen 1 721,81 valutaenheter.  
ÅRSAVSKR, LINAVSKR, VDEGRAVSKR.  
DB  
Beräknar avskrivningen enligt den geometrisk-degressiva metoden för en viss avskrivningstid.  
Den här avskrivningsformen använder Du när Du vill att avskrivningsvärdet ska vara störst i början av avskrivningen (i motsats till linjär avskrivning).  
Avskrivningsvärdet minskar med varje avskrivningsperiod med de avskrivningar som redan har dragits av från anskaffningsvärdet.  
Syntax  
DB( AV;RV;LL;P;MÅ)  
AV är tillgångens anskaffningsvärde.  
RV är tillgångens restvärde vid livslängdens slut.  
LL är livslängden uttryckt i antalet avskrivningsperioder.  
P är periodlängden.  
Du måste ange perioden i samma tidsenhet som livslängden.  
MÅ (valfritt) är antalet månader under första avskrivningsåret.  
Om inget annat anges används faktorn 12.  
Exempel  
Ett datorsystem med ett anskaffningsvärde på 25 000 valutaenheter ska skrivas av på tre år.  
Restvärdet ska vara 1 000 valutaenheter.  
En period utgörs av 30 dagar.  
DB( 25000;1000;36;1;6) = 1 075,00 valutaenheter  
Den geometriskt degressiva avskrivningen av datorsystemet är 1 075 valutaenheter.  
DEGAVSKR, VDEGRAVSKR, ÅRSAVSKR.  
IR  
Med den här funktionen kan du beräkna internräntan för en investering utan att ta hänsyn till kostnader eller intäkter.  
På det sättet kan du undersöka en investerings räntabilitet.  
Syntax  
IR( värden;gissning)  
värden är en matris eller cellreferens till celler vars innehåll motsvarar betalningarna.  
gissning (valfritt) är ett uppskattat värde på räntefotens startvärde.  
Exempel  
Om cellerna A1 - A4 antas innehålla värdena A1=-10000,A2=13500,A3=7600 respektive A4=1000, visas som resultat värdet 80,24%.  
NETNUVÄRDE, RÄNTA.  
RALÅN  
Med den här funktionen kan du beräkna hur höga räntorna blir vid konstanta amorteringar.  
Syntax  
RALÅN( Ränta; Period; Perioder_totalt; investering)  
Ränta definierar den periodiska räntesatsen.  
Period är antalet amorteringsperioder för beräkningen av räntorna.  
Perioder_totalt är det totala antalet amorteringsperioder.  
investering är investeringsbeloppet.  
Exempel  
Vid en kreditsumma på 120 000 valutaenheter med två års löptid och amortering månadsvis, med en räntesats på 12% efterfrågas hur höga räntorna är efter 1,5 år.  
RALÅN( 1;18;24;120000) = -30 000 valutaenheter.  
Summan av räntorna uppgår till 30 000 valutaenheter efter 1,5 år.  
Till finansfunktionerna del 2  
Till finansfunktionerna del 3  
Kategorin Information  
Här visas de funktioner som finns i kategorin Information med ett exempel.  
Funktionerna omfattar AKTUELL, CELL FORMEL, N, SAKNAS, VÄRDETYP, ÄREJTEXT, ÄRF, ÄRFEL, ÄRFORMEL, ÄRJÄMN_ADD, ÄRLOGISK, ÄRREF, ÄRSAKNAD, ÄRTAL, ÄRTEXT, ÄRTOM ÄRUDDA_ADD.  
De beskrivs nedan.  
Några exempel går bara att förklara med hjälp av en tabell.  
Använd i sådana fall följande tabell som utgångspunkt.  
C  
D  
2  
x-värde  
y-värde  
3  
-5  
-3  
4  
-2  
0  
5  
-1  
1  
6  
0  
3  
7  
2  
4  
8  
4  
6  
9  
6  
8  
AKTUELL  
Beräknar formelns aktuella värde, vid den position vid vilken denna funktion befinner sig.  
Syntax  
AKTUELL().  
Exempel  
Den här funktionen kan Du t ex använda tillsammans med cellformateringsfunktionen FORMATMALL när Du vill tilldela den aktuella cellen det aktuella värdet flr en ny formatering.  
=AKTUELL( )+FORMATMALL(Ny)  
1+2+AKTUELL() ger 6 (1+2=AKTUELL+AKTUELL=6)  
1+AKTUELL( )+2 ger 4 (1=AKTUELL+AKTUELL+2=4)  
FORMEL  
Funktionen visar formeln i en formelcell på ett godtyckligt ställe.  
Formeln i en formelcell returneras som sträng vid positionen Referens.  
Om det inte finns någon formelcell där eller om det överlämnade argumentet inte är någon referens sätts #Saknas.  
Syntax  
FORMEL()  
Exempel  
I cell A8 står värdet 23 som resultat av en formel.  
I cellen A1 kan Du t ex då utnyttja funktionen FORMEL för att visa formeln i cellen A8.  
=FORMEL( A8)  
ÄRREF  
Denna funktion kontrollerar om innehållet i en eller flera är en referens.  
Referenstyperna kontrolleras med avseende på såväl enskilda celler som cellområden.  
Syntax  
ÄRREF( värde)  
värde är det värde för vilket det ska kontrolleras om det rör sig om en referens.  
Exempel  
ÄRREF( C5) ger resultatet SANT.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRF  
Denna funktion ger resultatet SANT om den kontrollerade cellen ger ett felvärde som inte är lika med #Saknas.  
Denna informationsfunktion kan Du använda för att kontrollera förekomsten av felvärden i vissa celler.  
Syntax  
ÄRF( värde)  
värde är ett godtyckligt värde eller uttryck med vilket Du kontrollerar om det finns ett felvärde som inte är lika med #Saknas eller inte.  
Exempel  
ÄRF( C5) ger FALSKT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRFEL  
Till skillnad från ÄRF kontrollerar ÄRFEL om det överhuvudtaget finns felvärden i celler eller inte.  
ÄRFEL identifierar felvärdet #Saknas.  
Syntax  
ÄRFEL( värde)  
värde är ett godtyckligt uttryck, med vilket Du kontrollerar om det rör sig om ett felvärde eller inte.  
Exempel  
ÄRFEL( C8) ger FALSKT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRFORMEL  
Denna funktion kontrollerar om en cell innehåller en formel.  
Syntax  
ÄRFORMEL( referens)  
referens anger referensen till en cell, för vilken Du vill kontrollera om den innehåller en referens.  
Exempel  
ÄRFORMEL( D4) ger FALSKT som resultat.  
ÄRJÄMN_ADD  
Resultatet är SANT (1) om talet delat med 2 ger ett heltal som resultat, annars FALSKT (0).  
Syntax  
ÄRJÄMN_ADD( Tal)  
Tal: talet som ska kontrolleras.  
Exempel  
=ÄRJÄMN_ADD( 5) ger resultatet 0.  
ÄREJTEXT  
Kontrollerar om cellinnehållet är text eller siffror.  
Om cellinnehållet är text returneras resultatet FALSKT.  
Syntax  
ÄREJTEXT( värde)  
värde är ett värde eller ett uttryck för vilket Du vill kontrollera om det rör sig om en text, ett tal eller ett logiskt värde.  
Exempel  
ÄREJTEXT( D2) ger FALSKT som resultat.  
ÄREJTEXT( D9) ger SANT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRTOM  
Denna funktion ger resultatet SANT om cellreferensen är tom.  
Denna informationsfunktion använder Du för att kontrollera om innehållet i en cell är tomt.  
Syntax  
ÄRTOM( värde)  
värde är ett godtyckligt innehåll, som Du har angett i den cell som ska kontrolleras.  
Exempel  
ÄRTOM( D2) ger FALSKT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRLOGISK  
Den här funktionen ger SANT som resultat om det kontrollerade uttrycket har ett logiskt talformat.  
Du använder funktionen för att kontrollera förekomsten av de båda logiska värdena SANT och FALSKT i vissa celler.  
Syntax  
ÄRLOGISK( värde)  
värde är ett värde för vilket Du vill kontrollera om dess format motsvarar ett logiskt talformat.  
Exempel  
ÄRLOGISK( D5) ger FALSKT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRSAKNAD  
Kontrollerar om en cell innehåller felvärdet #Saknas (värdet är ej tillgängligt) och returnerar SANT om det kontrollerade felvärdet är #Saknas.  
Syntax  
ÄRSAKNAD( värde)  
värde är värdet eller ett uttryck som ska kontrolleras.  
Exempel  
ÄRTOM( D3) ger FALSKT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRTEXT  
Kontrollerar om cellinnehållet är text eller siffror.  
Returnerar SANT om cellinnehållet är en text.  
Syntax  
ÄRTEXT( värde)  
värde är ett värde, ett tal, ett logiskt värde eller ett felvärde för vilket kontrolleras om det är text eller tal.  
Exempel  
ÄRTEXT( C2) ger SANT som resultat.  
ÄRTEXT( C3) ger FALSKT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
ÄRUDDA_ADD  
Resultatet är SANT (1) om talet delat med 2 inte ger ett heltal som resultat, annars FALSKT (0).  
Syntax  
ÄRUDDA_ADD( Tal)  
Tal: talet som ska kontrolleras.  
Exempel  
=ÄRUDDA_ADD( 5) ger resultatet 1.  
ÄRTAL  
Denna funktion returnerar SANT om det kontrollerade värdet är ett tal.  
Syntax  
ÄRTAL( värde)  
värde är ett godtyckligt värde som ska kontrolleras för att se om det är ett tal eller en text.  
Exempel  
ÄRTAL( C3) ger SANT som resultat.  
ÄRTAL( C2) ger FALSKT som resultat.  
FELTYP, ÄRJÄMN, ÄRUDDA, VÄRDETYP.  
N  
Med denna funktion kan Du omvandla ett tal.  
Den här funktionen kan Du använda för att omvandla logiska värden till talvärdena 1 eller 0.  
Syntax  
N( värde)  
värde är ett värde som ska omvandlas till ett tal.  
Exempel  
N( SANT) returnerar 1  
N( FALSKT) returnerar 0  
N( #Saknas) returnerar 0  
T.  
SAKNAS  
Den här funktionen returnerar felvärdet #Saknas för en cell.  
Syntax  
SAKNAS()  
Exempel  
SAKNAS() omvandlar cellinnehållet till #Saknas.  
ÄRREF, ÄRF, ÄRFEL, ÄRFORMEL.  
ÄREJTEXT, ÄRTOM, ÄRLOG, ÄRSAKNAD, ÄRTEXT, ÄRTAL.  
VÄRDETYP  
Fastställer ett värdes datatyp.  
Syntax  
VÄRDETYP( värde)  
värde är ett visst värde för vilken datatypen ska fastställas. värde 1 = tal, värde 2 = text, värde 4 = logiskt värde, värde 8 = formel, värde 16 = felvärde.  
Exempel (se exempeltabell ovan)  
VÄRDETYP( C2) returnerar 2 som resultat.  
VÄRDETYP( D9) returnerar 1 som resultat.  
CELL  
Ger information om adress, formatering eller innehåll i en cell.  
Syntax  
CELL( infotyp; referens)  
infotyp är strängen som bestämmer informationstypen.  
Strängen är alltid på engelska och inte versalkänslig.  
info_typ  
Betydelse  
COL  
Returnerar numret på den refererade kolumnen.  
Cell( "COL";D2) returnerar 4.  
ROW  
Returnerar numret på den refererade raden.  
Cell( "ROW";D2) returnerar 2.  
SHEET  
Returnerar numret på den refererade tabellen.  
CELL( "Sheet";Tabell3.D2) returnerar 3.  
ADRESS  
Returnerar den absoluta adressen på den refererade tabellen.  
CELL( "ADDRESS";D2) returnerar $D$2.  
CELL( "ADDRESS";Tabell3.D2) returnerar $Tabell3.$D$2.  
CELL( "ADDRESS" ;'X:\dr\test.sxc'#$Tabell1.D2) returnerar 'file: / //X: / dr / test.sxc '#$Tabell1.$D$2.  
FILENAME  
Returnerar filnamn och tabellnamn på den refererade cellen.  
CELL( "FILENAME";D2) returnerar 'file: / //X: / dr / own.sxc '#$Tabell1 om formeln i det aktuella dokumentet X:\dr\own.sxc står i Tabell1.  
CELL( "FILENAME" ;'X:\dr\test.sxc'#$Tabell1.D2) returnerar 'file: / //X: / dr / test.sxc '#$Tabell1.  
COORD  
Returnerar den fullständiga celladressen i Lotus( TM )-beteckningssätt.  
CELL( "COORD"; D2) returnerar $A:$D$2.  
CELL( "COORD"; Tabell3.D2) returnerar $C:$D$2.  
CONTENTS  
Returnerar innehållet i den refererade cellen utan någon formatering.  
TYPE  
Returnerar typen av cellinnehåll.  
b = blank. tom cell  
l = label.  
Text, resultat av en formel i form av text  
v = value.  
Värde, resultat av en formel i form av tal  
WIDTH  
Returnerar bredden på den refererade kolumnen.  
Måttenheten är antalet nollor (0) som passar i kolumnen, i standardteckensnittet med standardstorlek.  
PREFIX  
Returnerar justeringen på den refererade cellen.  
'= vänsterjusterad eller marginaljusterad  
"= högerjusterad  
^ = centrerad  
\ = upprepande (inaktiv för närvarande)  
PROTECT  
Returnerar status för cellens cellskydd.  
1 = cell är skyddad  
0 = cell är inte skyddad  
FORMAT  
Returnerar en sträng som anger talformatet.  
, = tal med tusentalsavgränsare  
F = tal utan tusentalsavgränsare  
C = valutaformat  
S = exponentiell framställning, t.ex. 1.234+E56  
P = procenttal  
I de ovannämnda formaten anges antalet decimaler som tal efter decimaltecknen.  
Exempel:  
Talformatet #,##0.0 returnerar ,1 och talformatet 00.000% returnerar P3  
D1 = D-MMM-YY, D-MM-YY och liknande format  
D2 = DD-MM  
D3 = MM-YY  
D4 = DD-MM-YYYY HH:MM:SS  
D5 = MM-DD  
D6 = HH:MM:SS AM / PM  
D7 = HH:MM AM / PM  
D8 = HH:MM:SS  
D9 = HH:MM  
G = Alla andra format  
- (minus) i slutet = negativa tal formateras med färg  
() (parentespar) i slutet = det förekommer en inledande parentes i formatkod  
COLOR  
Returnerar 1 om negativa värden är formaterade med färg, annars 0.  
PARENTHESES  
Returnerar 1 om det finns en öppen parentes (i formatkoden, annars 0.  
referens (valfritt) är positionen för cellen som ska undersökas.  
Om referens är ett område, gäller cellen uppe till vänster i området.  
Om referens saknas, använder %PRODUCTNAME Calc positionen för cellen där den här formeln står.  
Microsoft Excel använder då referensen för cellen där markören står.  
Kategorin Logisk  
Här visas de funktioner som är tillgängliga i kategorin Logisk med ett exempel.  
Det rör sig om funktionerna FALSKT, ICKE, ELLER, OCH, SANT och OM.  
De beskrivs nedan.  
FALSKT  
Med det här kommandot bestämmer Du det logiska värdet för falskt.  
Två eller fler argument länkas med de logiska operatorerna OCH eller ELLER.  
Länken ger det logiska värdet FALSKT om argumentens innehåll kräver detta.  
Syntax  
FALSKT()  
Exempel  
Om A=SANT och B=FALSKT erhåller Du följande exempel:  
A OCH B returnerar FALSKT  
A ELLER B returnerar SANT  
SANT.  
ICKE  
Med den här funktionen kastas det logiska värdet om.  
Syntax  
ICKE (logiskt värde)  
Det logiska värdet är ett godtyckligt värde som ska kastas om.  
Exempel  
ICKE( A).  
A=SANT ger då A=FALSKT.  
ELLER, OCH.  
ELLER  
Returnerar SANT om minst ett argument är SANT.  
Om alla argument har värdet FALSKT returnerar den här funktionen FALSKT.  
Argumenten är antingen egna logiska uttryck (SANT, 1<5, 2+3=7, B8<10), som returnerar logiska värden, eller matriser (A1:C3), som innehåller logiska värden.  
Om ett argument som är angivet som en matris innehåller text eller tomma celler, ignoreras dessa värden.  
Formeln =ELLER( 0<C9:C16; FALSKT) returnerar t ex värdet SANT om matrisen (C9:C16) innehåller värden större än 0, varvid även celler med text eller tomma celler kan förekomma.  
Om det angivna området inte innehåller några logiska värden, returnerar ELLER felvärdet #Värde!.  
Syntax  
ELLER( logiskt värde 1; logiskt värde 2... logiskt värde 30)  
Logiskt värde 1; logiskt värde 2... logiskt värde 30 är villkor som ska undersökas.  
Varje villkor kan vara antingen SANT eller FALSKT.  
Om Du anger ett område som parameter, kopplas de enskilda logiska värdena i de celler som området innehåller ihop med operatorn ELLER.  
Resultatet är SANT om någon av cellerna i området har det logiska värdet SANT.  
Exempel  
Du ska undersöka posterna 12<11; 13>22 och 45=45 med avseende på deras logiska värden.  
ELLER( 12<11; 13>22; 45=45) returnerar SANT.  
ELLER( FALSKT;SANT) returnerar SANT.  
ICKE, OCH.  
OCH  
Returnerar SANT om alla argument har värdet SANT.  
Om ett argument har värdet FALSKT returnerar den här funktionen FALSKT.  
Argumenten är antingen egna logiska uttryck (SANT, 1<5, 2+3=7, B8<10), som returnerar logiska värden, eller matriser (A1:C3), som innehåller logiska värden.  
Om ett argument som är angivet som en matris innehåller text eller tomma celler, ignoreras dessa värden.  
Formeln =OCH( 0<C9:C16; C9:C16<10) returnerar t ex värdet SANT om matrisen (C9:C16) innehåller värden mellan 0 och 10, varvid även celler med text eller tomma celler kan förekomma.  
Om det angivna området inte innehåller några logiska värden, returnerar OCH felvärdet #VÄRDE!.  
Syntax  
OCH( logiskt värde 1; logiskt värde 2... logiskt värde 30)  
Logiskt värde 1; logiskt värde 2... logiskt värde 30 är villkor som ska undersökas.  
Varje villkor kan vara antingen SANT eller FALSKT.  
Om Du anger ett område som parameter, kopplas de enskilda logiska värdena i de celler som området innehåller ihop med operatorn OCH.  
Resultatet är SANT om alla celler i området har det logiska värdet SANT.  
Exempel  
Du ska undersöka posterna 12<13; 14>12 och 7<6 med avseende på deras logiska värden.  
OCH( 12<13; 14>12; 7<6) returnerar FALSKT.  
OCH (FALSKT;SANT) returnerar FALSKT.  
ICKE, ELLER.  
SANT  
Det logiska värdet SANT sätts.  
Den logiska funktionen SANT undersöker två argument och sätter det logiska värdet SANT om båda värdena stämmer överens.  
Syntax  
SANT()  
Exempel  
Om A=SANT och B=FALSKT erhåller Du följande exempel:  
A OCH B returnerar FALSKT  
A ELLER B returnerar SANT  
(ICKE) A OCH B returnerar SANT  
FALSKT  
OM  
Undersöker det logiska värdet på en Om-Så-koppling.  
Syntax  
OM( test; värde_om_sant; värde_om_falskt)  
test är ett godtyckligt värde eller uttryck som kan vara SANT eller FALSKT.  
värde_om_sant (valfritt) är funktionens resultat om det logiska testet ger resultatet SANT.  
värde_om_falskt (valfritt) är funktionens resultat om det logiska testet ger resultatet FALSKT.  
Exempel  
OM( A1>5;100 ;"för lågt") Om värdet i A1 är större än 5, införs i den aktuella cellen värdet 100, annars införs texten för lågt.  
FALSKT, ICKE, ELLER, OCH, SANT.  
Kategori Matematik  
Du får även ett exempel.  
Hur Du använder Funktionsautopiloten beskrivs får Du reda på via menyn Infoga - Funktion.  
Du har tillgång till följande funktioner:  
ABS, ANTAL.OM, ANTAL.TOMMA, ARCCOS, ARCCOSH, ARCCOT, ARCCOTH, ARCSIN, ARCSINH, ARCTAN, ARCTAN2, ARCTANH, AVKORTA, AVRUNDA, AVRUNDA.NEDÅT, AVRUNDA.UPPÅT, COS, COSH, COT, COTH, DELSUMMA, EXP, FAKULTET, GRADER, HELTAL, JÄMN, KOMBIN, KOMBIN2, KVADRATSUMMA, KVOT, LN, LOG, LOG10, MAVRUNDA, MGM, MGM_ADD, MULTINOMIAL, OMRÄKNA, PI, PRODUKT, RADIANER, REST, ROT, ROTPI, RUNDA.NER, RUNDA.UPP, SERIESUMMA, SIN, SINH, SGD, SGD_ADD, SLUMP, SLUMP.MELLAN, SUMMA, SUMMA.OM, TAN, TANH, TECKEN, UDDA, UPPHÖJT.TILL, ÄRJÄMN, ÄRUDDA,.  
En del funktioner avser tabellfunktioner.  
I dessa fall används följande tabell som utgångspunkt.  
A  
B  
C  
D  
E  
1  
167,56  
351,10  
57,25  
17,95  
870,29  
2  
479,01  
269,99  
86,30  
351,10  
3  
12,60  
22,50  
4  
AVRUNDA.NEDÅT  
Med den här funktionen avrundar Du ett tal nedåt till det antal decimaler som Du själv har definierat.  
Syntax:  
AVRUNDA.NEDÅT( tal; antal)  
tal är det tal som ska avrundas nedåt.  
antal (valfritt) är det antal decimaler som talet ska avrundas till.  
Om parametern antal är negativ, så sker avrundningen till siffror framför kommatecknet.  
Exempel:  
Om Du anger värdet 567,567 och skriver 2 i fältet antal blir resultatet 567,56.  
AVRUNDA.UPPÅT, HELTAL, AVKORTA, RUNDA.UPP, REST, AVRUNDA, RUNDA.NER  
ABS  
Här kan Du beräkna absolutvärdet för ett tal.  
Syntax:  
ABS( tal)  
tal är det värde vars absolutvärde ska beräknas.  
Exempel:  
Om Du anger värdet -56 blir absolutvärdet 56.  
Om Du anger värdet 56 blir absolutvärdet 56.  
TECKEN  
ANTAL.TOMMA  
Om Du vill ta reda hur många celler som inte har något innehåll, anger Du cellreferenserna åtskilda med kolon i textfältet område.  
Syntax:  
ANTAL.TOMMA( område)  
område är området där de tomma cellerna räknas.  
Exempel:  
Om Du anger = ANTAL.TOMMA (A1:C3) i ett tomt cellområde blir resultatet 9.  
ANTAL.OM  
ARCCOS  
Arcuscosinus beräknas utifrån det tal som du har angett i textfältet tal.  
Syntax:  
ARCCOS( tal)  
tal är det värde vars arcuscosinusvärde ska beräknas.  
Exempel:  
Arcuscosinus för -1 ger värdet 3,14.  
Arcuscosinus för 0 ger värdet 1,57.  
Arcuscosinus för 1 ger värdet 0.  
ARCSIN, ARCTAN, ARCCOT, COS  
ARCCOSH  
Ur det tal som Du anger i textfältet tal beräknas dess inversa hyperboliska cosinus.  
Syntax:  
ARCCOSH( tal)  
tal är värdet vars inversa hyperboliska cosinus ska beräknas.  
Exempel:  
Den inversa hyperboliska cosinus för 1 ger värdet 0.  
Den inversa hyperboliska cosinus för 15 ger värdet 3,4.  
Den inversa hyperboliska cosinus för 30 ger värdet 4,09.  
ARCSINH, ARCTANH, ARCCOTH, COSH  
ARCCOT  
Ur det tal som Du anger i textfältet tal beräknas arcuscotangens.  
Syntax:  
ARCCOT( tal)  
tal är värdet vars arcuscotangens ska beräknas.  
Exempel:  
Arcuscotangens för -1 ger värdet 2,36.  
Arcuscotangens för 0 ger värdet 1,57.  
Arcuscotangens för 1 ger värdet 0,79.  
ARCTAN, ARCSIN, ARCCOS, COT  
ARCCOTH  
Ur det tal som Du anger i textfältet tal beräknas dess inversa hyperboliska cotangens.  
Syntax:  
ARCCOTH( tal)  
tal är värdet vars inversa hyperboliska cotangens ska beräknas.  
Exempel:  
Den inversa hyperboliska cotangens för 1,1 ger värdet 1,52.  
Den inversa hyperboliska cotangens för 45 ger värdet 0,02.  
Den inversa hyperboliska cotangens för 90 ger värdet 0,01.  
ARCTANH, ARCSINH, ARCCOSH, COTH  
ARCSIN  
Ur det tal som Du anger i textfältet tal beräknas arcussinus.  
Syntax:  
ARCSIN( tal)  
tal är värdet vars arcussinusvärde ska beräknas.  
Exempel:  
Arcussinus för -1 ger värdet -1,57.  
Arcussinus för 0 ger värdet 0.  
Arcussinus för 1 ger värdet 1,57.  
ARCCOS, ARCTAN, ARCCOT, SIN  
ARCSINH  
Ur det tal som Du anger i textfältet tal beräknas dess inversa hyperboliska sinus.  
Syntax:  
ARCSINH( tal)  
tal är värdet vars inversa hyperboliska sinus ska beräknas.  
Exempel:  
Den inversa hyperboliska sinus för -90 ger värdet -5,19.  
Den inversa hyperboliska sinus för 0 ger värdet 0.  
Den inversa hyperboliska sinus för 90 ger värdet 5,19.  
ARCCOSH, ARCTANH, ARCCOTH, SINH  
ARCTAN  
Arcustangens beräknas ur det tal som Du anger i textfältet tal.  
Syntax:  
ARCTAN( tal)  
tal är det värde vars arcustangensvärde Du ska beräkna.  
Exempel:  
Arcustangens för -1 ger värdet -0,79.  
Arcustangens för 0 ger värdet 0.  
Arcustangens för 45 ger värdet 1,55.  
ARCSIN, ARCCOS, ARCCOT, TAN, ARCTAN2  
ARCTAN2  
Om Du vill ha arcustangens i koordinatvisning, anger Du värdet för x-koordinaten i textfältet tal_x och värdet för y-koordinaten i textfältet tal_y.  
Syntax:  
ARCTAN2( tal_x; tal_y)  
tal_x är värdet för x-koordinaten.  
tal_y är värdet för y-koordinaten.  
Exempel:  
Om Du anger värdet 45 för x-koordinaten och värdet 90 för y-koordinaten blir arcustangens 1,11.  
Om Du anger värdet -1 för x-koordinaten och värdet 0 för y-koordinaten blir arcustangens 3,14.  
ARCTAN, ARCTANH, PI, TAN  
ARCTANH  
Ur det tal som Du anger i textfältet tal beräknas dess inversa hyperboliska tangens.  
Syntax:  
ARCTANH( tal)  
tal är värdet vars inversa hyperboliska tangens ska beräknas.  
Exempel:  
Den inversa hyperboliska tangens för 0,99 ger värdet 2,65.  
Den inversa hyperboliska tangens för 0 ger värdet 0.  
Den inversa hyperboliska tangens för -0,95 ger värdet -1,83.  
ARCCOTH, ARCSINH, ARCCOSH, TANH  
AVRUNDA.UPPÅT  
Med den här funktionen kan Du avrunda ett tal uppåt till antal decimaler som Du själv har angett.  
Syntax:  
AVRUNDA.UPPÅT( tal; antal)  
tal är talet som ska avrundas uppåt.  
antal (valfritt) är antalet decimaler som talet ska avrundas till.  
Exempel:  
Om Du anger värdet 123,343 och skriver 2 i fältet antal blir resultatet 123,35.  
AVRUNDA.NEDÅT, HELTAL, AVKORTA, RUNDA.UPP, REST, AVRUNDA, RUNDA.NER  
COS  
Cosinus för en vinkel beräknas ur det tal som Du anger i textfältet tal.  
Syntax:  
COS( tal)  
tal är det värde vars cosinus ska beräknas.  
Exempel:  
Vinkeln 6,28 (2pi) mätt i bågmåttet ger cosinus på 1.  
Vinkeln 3,14 (pi) mätt i bågmåttet ger cosinus på -1.  
Vinkeln 1,57 (pi / 2) mätt i bågmåttet ger cosinus på 0.  
SIN, TAN, COT, PI, ARCCOS  
COSH  
Ur det tal som Du anger i textfältet tal beräknas den hyperboliska cosinus för en vinkel.  
Syntax:  
COSH( tal)  
tal är värdet vars hyperboliska cosinus ska beräknas.  
Exempel:  
Om Du anger värdet -5 blir den hyperboliska cosinus 74,21.  
Om Du anger värdet 0 blir den hyperboliska cosinus 1.  
Om Du anger värdet 90 blir den hyperboliska cosinus 6,10E038.  
SINH, TANH, COTH, ARCCOSH  
COT  
Ur det tal som Du anger i textfältet beräknas cotangens för en vinkel.  
Syntax:  
COT( tal)  
tal är det värde vars cotangens Du ska beräkna.  
Exempel:  
Vinkeln -45 mätt i bågmåttet ger cotangens på -0,62.  
Vinkeln 90 mätt i bågmåttet ger cotangens på -0,5.  
SIN, COS, TAN, PI, ARCCOT  
COTH  
Ur det tal som Du anger i textfältet tal beräknas den hyperboliska cotangens för en vinkel.  
Syntax:  
COTH( tal)  
tal är värdet vars hyperboliska cotangens ska beräknas.  
Exempel:  
Om Du anger värdet 90 blir den hyperboliska cotangens 1.  
Om Du anger värdet 45 blir den hyperboliska cotangens 1.  
Om Du anger värdet -45 blir den hyperboliska cotangens -1.  
TANH, SINH, COSH, ARCCOTH  
GRADER  
Ur det bågmått (radianer) som Du anger i textfältet tal beräknas gradtalet för vinkeln.  
Syntax:  
GRADER( tal)  
tal är värdet vars gradtal ska beräknas.  
Exempel:  
Ur det inmatade värdet 0,1 beräknas graderna till 5,73 för vinkeln.  
Ur det inmatade värdet 1,5708 beräknas graderna till 90 för vinkeln.  
Ur det inmatade värdet -0,7854 beräknas graderna till -45 för vinkeln.  
RADIANER, PI  
EXP  
Ur det värde som Du anger i textfältet beräknas exponenten för basen e.  
Syntax:  
EXP( tal)  
tal är exponenten till basen e.  
Exempel:  
Exponenten till basen e för värdet -4 ger som resultat 0,02.  
Exponenten till basen e för värdet 0,5 ger som resultat 1,65.  
Exponenten till basen e för värdet 1 ger som resultat 2,72.  
LN, LOG, UPPHÖJT.TILL  
FAKULTET  
Ur det värde som Du anger i textfältet tal beräknas fakulteten.  
Syntax:  
FAKULTET( tal)  
tal är det värde vars fakultet Du ska beräkna.  
Exempel:  
Fakulteten för talet 0 är 1.  
Fakulteten för värdet 3 är 6.  
Fakulteten för värdet 10 är 3628880.  
PRODUKT  
HELTAL  
Det tal som Du anger i textfältet avrundas nedåt till närmaste mindre heltal.  
Syntax:  
HELTAL( tal)  
tal är talet som ska avrundas nedåt till närmast mindre heltal.  
Exempel:  
Om Du anger talet -0,1 blir resultatet -1.  
Om Du anger talet 23,74 blir resultatet 23.  
AVKORTA, RUNDA.UPP, REST, AVRUNDA, RUNDA.NER  
JÄMN  
Det tal som Du anger i textfältet tal avrundas uppåt till närmaste jämna heltal.  
Syntax:  
JÄMN( tal)  
tal är talet som ska avrundas uppåt till närmaste jämna heltal.  
Exempel:  
Om Du anger talet 0,01 blir resultatet 2.  
Om Du anger talet -2,1 blir resultatet -4.  
Om Du anger talet 17,9 blir resultatet 18.  
HELTAL, ÄRJÄMN, ÄRUDDA, AVKORTA, RUNDA.UPP, AVRUNDA, UDDA, RUNDA.NER  
SGD  
Om Du ur olika tal vill bestämma deras största gemensamma nämnare, så anger Du de tal som ska jämföras i textfälten heltal.  
Syntax:  
SGD( heltal 1 till 30)  
Heltal 1 till 30 är upp till 30 heltal vars största gemensamma nämnare ska beräknas.  
Exempel:  
Om Du matar in talen 512, 1024 och 2000 i textfälten heltal 1, 2 och 3, visas 16 som resultat.  
MGM  
SGD_ADD  
Resultatet är den största gemensamma täljaren i en lista med tal.  
Syntax  
SGD_ADD( Tal)  
Tal: en lista med upp till 30 tal.  
Exempel  
=SGD_ADD( 5;15;25) ger resultatet 5.  
ÄRJÄMN  
Om Du vill kontrollera om ett värde hör till de jämna talen, skriver Du in det i textfältet värde.  
E jämnt värde resulterar i svaret SANT, och ett udda i svaret FALSKT.  
Syntax:  
ÄRJÄMN( värde)  
värde är värdet som ska kontrolleras.  
Exempel:  
När Du har angett värdet 642 visas SANT som resultat.  
Om Du anger värdet -4 visas SANT som resultat.  
Om Du anger värdet 7,6 visas FALSKT som resultat.  
JÄMN, ÄRUDDA, UDDA  
ÄRUDDA  
Om Du vill kontrollera om ett värde hör till de udda talen, skriver Du in det i textfältet värde.  
För ett udda värde visas svaret SANT, och för ett jämnt visas svaret FALSKT.  
Syntax:  
ÄRUDDA( värde)  
värde är värdet som ska kontrolleras.  
Exempel:  
Om Du anger värdet 642 visas FALSKT som resultat.  
Om Du anger värdet -4 visas FALSKT som resultat.  
Om Du anger värdet 7,6 visas SANT som resultat.  
JÄMN, ÄRJÄMN, UDDA  
MGM  
Om Du ur olika tal vill bestämma deras minsta gemensamma multipel, så anger Du i textfälten heltal de tal som ska jämföras.  
Syntax:  
MGM( heltal 1 till 30)  
Heltal 1 till 30 är upp till 30 heltal vars minsta gemensamma multipel ska beräknas.  
Exempel:  
Om Du anger talen 512, 1024 och 2000 i textfälten heltal 1, 2 och 3, visas 128000 som resultat.  
SGD  
MGM_ADD  
Resultatet är den minsta gemesamma multipeln i en lista med tal.  
Syntax  
MGM_ADD( Tal)  
Tal: en lista med upp till 30 tal.  
Exempel  
=MGM_ADD( 5;15;25) ger resultatet 75.  
KOMBIN  
Här kan Du beräkna antalet elementkombinationer utan upprepning.  
Syntax:  
KOMBIN( antal_1; antal_2)  
antal_1 är det totala antalet element.  
antal_2 är det valda antalet element.  
Exempel:  
Om Du anger talet 2 i textfälten antal_1 och antal_2 visas 1 som resultat.  
KOMBIN2, BINOMFÖRD, FAKULTET, HYPGEOMFÖRD, KRITBINOM, NEGBINOMFÖRD, PERMUT  
KOMBIN2  
Här kan Du beräkna antalet kombinationer av element med upprepning.  
Syntax:  
KOMBIN2( antal_1; antal_2)  
antal_1 är det totala antalet element.  
antal_2 är det utvalda antalet element.  
Exempel:  
Om Du skriver talet 2 i textfälten antal_1 och antal_2 visas 3 som resultat.  
KOMBIN, BINOMFÖRD, FAKULTET, HYPGEOMFÖRD, KRITBINOM, NEGBINOMFÖRD, PERMUT2  
AVKORTA  
Om Du vill avkorta ett tal till det antal decimaler som anges i textfältet antal, så skriver Du in detta tal i textfältet tal.  
När du anger antalet decimaler bör du kontrollera antalet decimaler som du har angett under Verktyg - Alternativ - Tabelldokument - Beräkna i fältet Antal decimaler.  
Ändra detta värde så att det motsvarar det önskade antalet decimaler.  
Syntax:  
AVKORTA( tal; antal)  
tal är talet vars decimaler ska avkortas.  
antal är antalet decimaler som inte ska avkortas.  
Exempel:  
Om Du skriver talet 34,5678 och antalet 1 visas 34,5 som resultat.  
Om Du skriver talet -15,769 och antalet 2, visas -15,77 som resultat.  
HELTAL, RUNDA.UPP, REST, AVRUNDA, RUNDA.NER  
LN  
Ur det värde som Du anger i textfältet beräknas den naturliga logaritmen för basen e.  
Syntax:  
LN( tal)  
tal är värdet vars naturliga logaritm ska beräknas.  
Exempel:  
Den naturliga logaritmen för basen e för värdet 3 ger som resultat 1,1.  
Den naturliga logaritmen för basen e för värdet 13 ger som resultat 2,56.  
Den naturliga logaritmen för basen e för värdet 1000 ger som resultat 6,91.  
EXP, LOG, LOG10  
LOG  
Ur det värde som Du anger i textfältet tal beräknas logaritmen för en valfri bas.  
Syntax:  
LOG( tal; bas)  
tal är det värde vars logaritm Du ska beräkna.  
bas är basen för logaritmberäkningen.  
Exempel:  
Logaritmen för talet 10 och basen 3 ger som resultat 2,1.  
Logaritmen för talet 2,1 och basen 7 ger som resultat 0,38.  
Logaritmen för talet 0,75 och basen 7,5 ger som resultat -0,14.  
EXP, LN, LOG10  
LOG10  
Ur det värde som Du anger i textfältet beräknas logaritmen för basen 10.  
Syntax:  
LOG10( tal)  
tal är värdet vars logaritm för basen 10 ska beräknas.  
Exempel:  
Logaritmen för basen 10 för värdet 3 ger som resultat 0,48.  
Logaritmen för basen 10 för värdet 10 ger som resultat 1.  
Logaritmen för basen 10 för värdet 0,02 ger som resultat -1,7.  
EXP, LN, LOG  
RUNDA.UPP  
Avrundar ett tal uppåt till närmaste signifikanta multipel.  
Syntax:  
RUNDA.UPP( tal, signifikans;läge)  
tal är talet som ska avrundas uppåt.  
signifikans är talet till vars multipel värdet ska avrundas uppåt.  
läge är ett valfritt värde.  
Om Du anger värdet och det ej är lika med noll, så avrundas talet beloppsmässigt uppåt vid negativt tal och signifikans.  
Observera att denna uppgift kan gå förlorad om Du exporterar till MS Excel eftersom Excel inte hanterar någon tredje parameter för funktioner.  
Om de båda parametrarna tal och signifikans är negativa och om värdet för läge är lika med noll eller inte har angetts, så är resultaten i %PRODUCTNAME Calc och i Excel olika efter export.  
Exempel:  
Om du skriver talet 3,4 och signifikansen 1 visas 4 som resultat.  
Om du matar in talet -6 och signifikansen -5 visas -5 som resultat.  
Om du skriver talet -0,6 och signifikansen -0,4 visas -0,4 som resultat.  
AVRUNDA.NEDÅT, AVRUNDA.UPPÅT, HELTAL, JÄMN, AVKORTA, AVRUNDA, UDDA, RUNDA.NER  
PI  
Här visas värdet pi (3,14...).  
Syntax:  
PI()  
Exempel:  
Pi motsvarar det avrundade värdet 3,14...  
SIN, COS  
MULTINOMIAL  
Returnerar fakulteten av en summa av argument delad med produkten av fakulteter av argument.  
Syntax  
MULTINOMIAL( Tal)  
Tal: en lista med upp till 30 tal.  
Exempel  
=MULTINOMIAL( F11:H11) ger resultatet 1260, om värdena 2, 3 och 4 står i F11 till H11.  
Det motsvarar formeln =( 2 !+3 !+4!) / 2!*3!*4!.  
UPPHÖJT.TILL  
Här kan Du upphöja ett tal till en exponent.  
Syntax:  
UPPHÖJT.TILL( bas; potens) eller bas ^ potens  
bas är talet som ska upphöjas.  
potens är exponenten som basen ska upphöjas till.  
Exempel:  
Om Du anger basen 3 och potensen -2 visas 0,11 som resultat.  
Om Du anger basen -3 och potensen -2 visas 0,11 som resultat.  
Om Du anger basen -3 och potensen 2 visas 9 som resultat.  
EXP, PRODUKT, ROT  
SERIESUMMA  
Ger en summa av potenser av tal x enligt följande formel som resultat:  
SERIESUMMA( x;n;m;Koefficienter) = Koefficient1xn + Koefficient2x(n+m) + Koefficient3x(n+2m) +... + Koefficientix(n+(i-1)m)  
Syntax  
x: talet som oberoende variabel  
n; initialpotens  
m: inkrementet  
Koefficienter: en serie koefficienter.  
Potensserien utökas med en del för varje koefficient.  
Exempel  
=SERIESUMMA( C12;D12;E12;F12:I12) ger resultatet 0,707103 (cosinus av PI / 4 radian eller 45 grader) om följande gäller: i C12 står =PI() / 4, i D12 står 0, i E12 står 2, i F12 står 1, i G12 står -1 / FAKULTET(2), i H12 står 1 / FAKULTET(4), i I12 står -1 / FAKULTET(6).  
PRODUKT  
Om Du ur flera tal vill beräkna deras produkt (multiplikation av argumenten), så skriver Du talen i textfälten tal.  
Syntax:  
PRODUKT( tal 1 till tal 30)  
tal 1 till tal 30 är upp till 30 argument vars produkt Du ska beräkna.  
Exempel:  
Om Du skriver talen 2, 3 och 4 i textfälten tal 1, 2 och 3, visas 24 som resultat.  
FAKULTET, SUMMA, PRODUKTSUMMA  
KVADRATSUMMA  
Om Du vill beräkna en kvadratsumma för några tal (summering av argumentens kvadrater), så skriver Du talen i textfälten.  
Syntax:  
KVADRATSUMMA( tal 1 till 30)  
tal 1 till tal 30 är upp till 30 argument vars kvadratsumma ska beräknas.  
Exempel:  
Om Du skriver talen 2, 3 och 4 i textfälten tal 1, 2 och 3, visas 29 som resultat.  
SUMMA, PRODUKTSUMMA  
KVOT  
Resultatet är heltalsresultatet av en division.  
Syntax  
KVOT( täljare;nämnare)  
Exempel  
=KVOT( 11;3) ger resultatet 3.  
Resten av 2 bortfaller.  
RADIANER  
Ur det gradtal som anges i textfältet beräknas bågmåttet (radianer).  
Syntax:  
RADIANER( tal)  
tal är vinkeln i grader.  
Exempel:  
Ur det angivna gradtalet 5,73 beräknas bågmåttet 0,1 för vinkeln.  
Ur det angivna gradtalet 90 beräknas bågmåttet 1,57 för vinkeln.  
Ur det angivna gradtalet -45 beräknas bågmåttet -0,79 för vinkeln.  
GRADER, PI  
REST  
Här kan Du beräkna restvärdet vid division med ett heltal.  
Syntax:  
REST( dividend; divisor)  
Dividend är det tal som ska delas.  
Divisor är talet som det ska divideras med.  
Exempel:  
Värdet 17 i fältet Dividend delas med divisorn -1,4.  
Som restvärde visas -1,2.  
Värdet -13 i fältet Dividend delas med divisorn -3,4.  
Som restvärde visas -2,8.  
Värdet 2987 i fältet Dividend delas med divisorn 362.  
Som restvärde visas 91.  
AVRUNDA.NEDÅT, AVRUNDA.UPPÅT, HELTAL, AVKORTA, AVRUNDA  
AVRUNDA  
Om du vill avrunda ett tal till ett visst antal decimaler enligt matematiskt giltiga kriterier, så anger du värdet i textfältet tal och det antal decimaler som talet ska avrundas till.  
Syntax:  
AVRUNDA( tal; antal)  
tal är talet som ska avrundas.  
antal (valfritt) är det antal decimaler som talet ska avrundas till.  
Om parametern antal är negativ, så sker avrundningen till siffror framför kommatecknet.  
Exempel:  
Om Du skriver talet 17,546 i fältet tal och antalet 1, visas 17,5 som resultat.  
Om Du skriver talet -32,483 i fältet tal och antalet 3 visas -32,48 som resultat.  
AVRUNDA.NEDÅT, AVRUNDA.UPPÅT, HELTAL, AVKORTA, RUNDA.UPP, REST, RUNDA.NER  
SIN  
Ur det tal som Du anger i textfältet tal beräknas sinus för en vinkel.  
Syntax:  
SIN( tal)  
tal är vinkeln i radianer (bågmått).  
Exempel:  
Vinkeln 3,14 (pi) mätt i radianer ger sinus på 0.  
Vinkeln 1,57 (pi / 2) mätt i radianer ger sinus på 1.  
Vinkeln 0,79 (pi / 4) mätt i radianer ger sinus på 0,71.  
COS, COT, TAN, PI, ARCSIN  
SINH  
Ur det tal som anger i textfältet tal beräknas den hyperboliska sinus för en vinkel.  
Syntax:  
SINH( tal)  
tal är talet vars hyperboliska sinus ska beräknas.  
Exempel:  
Om du anger värdet -5 blir den hyperboliska sinus -74,2.  
Om Du anger värdet 0 blir den hyperboliska sinus 0.  
Om Du anger värdet 90 ger den hyperboliska sinus 6,10E038.  
COSH, TANH, COTH, ARCSINH  
SUMMA  
Om Du vill beräkna argumentens summa ur flera tal, så skriver Du talen i textfälten tal.  
Syntax:  
SUMMA( tal 1; tal 2;...; tal 30)  
tal 1 till tal 30 är upp till 30 argument vars summa ska beräknas.  
Exempel:  
Om Du anger talen 2, 3 och 4 i textfälten tal 1, 2 och 3, visas 9 som resultat.  
SUMMA( A1;A3;B5) beräknar summan för de tre cellerna.  
SUMMA( A1:E10) beräknar summan för alla celler i cellområdet A1 till E10.  
Med funktionen SUMMA() kan Du använda villkor som är länkade med OCH tillsammans på följande sätt:  
Anta att Du har registrerat Dina räkningar i en tabell.  
I kolumn A står räkningarnas datum och i kolumn B beloppen.  
Du söker en formel med vilken Du kan summera enbart beloppen för en vissa månad, t ex beloppen för tidsintervallet >=1 januari 1999 till <1 februari 1999.  
Området med datum kan vara A1:A40 och området med de belopp som ska summeras kan vara B1:B40.  
I C1 står startdatumet för de räkningar som ska tas med, 1 januari 1999, och i C2 det datum som inte ska tas med, dvs den 1 februari 1999.  
Ange följande formel som matrisformel:  
=SUMMA( (A1:A40>=C1)*(A1:A40<C2)*B1:B40)  
Om Du vill ange den som matrisformel måste Du trycka ned Skift + Kommando Ctrl +Retur i stället för att bara avsluta med Retur.  
Formeln visas sedan i formellisten inom klammerparentes:  
{=SUMMA((A1:A40>=C1)*(A1:A40<C2)*B1:B40)}  
Formeln bygger på att resultatet av en jämförelse är 1 om kriteriet uppfylls och 0 om det inte uppfylls.  
De enskilda jämförelseresultaten behandlas däremot som matris och används i matrismultiplikationer och till slut summeras de enskilda värdena i resultatmatrisen.  
På detta sätt kan Du t ex även använda funktionen SUMMA() som ANTAL.OM() med flera kriterier.  
ANTAL, ANTALV, MEDEL, PRODUKT  
SUMMA.OM  
Om argumentens summa ska beräknas enbart om vissa villkor är uppfyllda, så anger Du område, kriterier och, om Du vill, summaområde.  
Den här funktionen kan Du använda för att genomsöka ett område efter ett visst värde.  
Syntax:  
SUMMA.OM( område; kriterier; summaområde)  
område är området som kriterierna ska tillämpas på.  
kriterier är den cell där sökkriteriet har angetts, eller själva sökkriteriet.  
summaområde är det område ur vilket värdena summeras.  
Om Du inte anger den här parametern, så summeras de värden som hittats i området.  
Exempel:  
Kriteriet 351,10 ska summeras ur området A1:E4 i exempeltabellen.  
Ange A1:E4 i textfältet område och som kriterium 351,10 eller B1.  
702,2 visas som resultat eftersom alla celler med innehållet 351,10 summeras.  
Tänk Dig att Du har en tabell i vilken Du hanterar Dina dagliga utgifter.  
I kolumn A (område) anges en kategori för varje enskilt kvitto, t ex "livsmedel", "tidskrifter "eller "reskostnader", och i kolumn B (summaområde) anges alltid beloppet för motsvarande kvitton.  
Formeln är: =SUMMA.OM( A1:A100 ;"livsmedel";B1:B100).  
Ytterligare ett exempel finns vid SUMMA().  
SUMMA, ANTAL.OM  
TAN  
Tangens för en vinkel beräknas ur det tal som Du har angett i textfältet.  
Syntax:  
TAN( tal)  
tal är vinkeln i radianer (bågmått).  
Exempel:  
Vinkeln 3,14 (pi) mätt i radianer ger tangens på 0.  
Vinkeln 0,79 (pi / 4) mätt i radianer ger tangens på 1,01.  
Vinkeln 0,39 (pi / 8) mätt i radianer ger tangens på 0,41.  
SIN, COS, COT, PI, ARCTAN  
TANH  
Ur det tal som Du anger i textfältet tal beräknas den hyperboliska tangens för en vinkel.  
Syntax:  
TANH( tal)  
tal är talet vars hyperboliska tangens ska beräknas.  
Exempel:  
Om Du anger värdet -5 blir den hyperboliska tangens -1.  
Om Du anger värdet 45 blir den hyperboliska tangens 1.  
Om Du anger värdet 90 blir den hyperboliska tangens 1.  
COTH, SINH, COSH, ARCTANH  
DELSUMMA  
Den här funktionen beräknar delresultat.  
Om området redan innehåller andra delresultat, används de inte i de fortsatta beräkningarna.  
Den här funktionen passar bra om du använder AutoFilter och bara vill ta hänsyn till de filtrerade dataposterna.  
Syntax:  
DELSUMMA( funktion; område)  
funktion är ett tal som står en av de följande funktionerna:  
Funktionsindex  
Funktion  
1  
MEDEL  
2  
ANTAL  
3  
ANTALV  
4  
MAX  
5  
MIN  
6  
PRODUKT  
7  
STDAV  
8  
STDAVP  
9  
SUMMA  
10  
VARIANS  
11  
VARIANSP  
område är det område vars celler ska inkluderas.  
Exempel:  
Antag att Du har en tabell i cellområdet A1:B5 med städer i kolumn A och tillhörande tal i kolumn B.  
Du har använt ett AutoFilter för att t ex bara visa de rader där staden är = "Hamburg".  
Följande formel skulle då passa väl:  
=DELSUMMA( 9; B2:B5)  
OMRÄKNA  
Med den här funktionen räknar du om ett valutavärde (t.ex. österrikiska schilling) till euro och omvänt.  
Omräkningsfaktorerna är sparade i filen calc.xml som finns i katalogen {installpath} / share / config / registry / instance / org / openoffice / Office.  
Syntax:  
OMRÄKNA( Värde ;"text" ;"text")  
värde är det valutabelopp som ska räknas om.  
text är beteckningen för den aktuella valutan och euron i ordningsföljden "från enhet" "till enhet ".  
Ange texten inom citattecken och ta hänsyn till versaler och gemener (t ex "EUR").  
Exempel:  
=OMRÄKNA( 100 ;"ATS" ;"EUR")  
=OMRÄKNA( 100 ;"EUR" ;"DEM")  
I tabellen hittar du valutabeteckningarna och de fixerade växelkurserna för euron som Europeiska kommissionen har fastlagt.  
Beräkningsbasen är 1 euro.  
Mer information hittar du på http: / /europa.eu.int / eurobirth / rates.html.  
"EUR"  
"ATS"  
13.7603  
Österrikiska schilling  
"EUR"  
"BEF"  
40.3399  
Belgiska franc  
"EUR"  
"DEM"  
1.95583  
Tyska mark  
"EUR"  
"ESP"  
166.386  
Spanska pesetas  
"EUR"  
"FIM"  
5.94573  
Finska mark  
"EUR"  
"FRF"  
6.55957  
Franska franc  
"EUR"  
"IEP"  
0.787564  
Irländska pund  
"EUR"  
"ITL"  
1936.27  
Italienska lire  
"EUR"  
"LUF"  
40.3399  
Luxemburgska franc  
"EUR"  
"NLG"  
2.20371  
Nederländska gulden  
"EUR"  
"PTE"  
200.482  
Portugisiska escudo  
"EUR"  
"GRD"  
340.750  
Grekisk drakma  
UDDA  
Det tal som Du anger i textfältet tal avrundas uppåt till närmaste udda heltal.  
Syntax:  
UDDA( tal)  
tal är det tal som ska avrundas uppåt.  
Exempel:  
Om Du anger talet 1,01 visas 3 som resultat.  
Om Du anger talet -3,01 visas -5 som resultat.  
Om Du anger talet 17,9 visas 19 som resultat.  
HELTAL, JÄMN, ÄRJÄMN, ÄRUDDA, AVKORTA, RUNDA.UPP, AVRUNDA, RUNDA.NER  
RUNDA.NER  
När Du vill avrunda ett tal till närmaste multipel av signifikansen, anger Du talet i textfältet tal och den önskade signifikansen i textfältet signifikans.  
Syntax:  
RUNDA.NER( tal, signifikans;läge)  
tal är det tal som ska avrundas nedåt.  
signifikans är det tal till vars multipel värdet ska avrundas nedåt.  
läge är ett valfritt värde.  
Om Du anger värdet och det ej är lika med noll, så avrundas talet beloppsmässigt uppåt vid negativt tal och signifikans.  
Det kan hända att detta värde ignoreras om Du exporterar till MS Excel eftersom Excel inte hanterar någon tredje parameter för funktioner.  
Om de båda parametrarna tal och signifikans är negativa och om värdet för läge är lika med noll eller inte har angetts, så är resultaten i %PRODUCTNAME Calc och i Excel olika efter export.  
Exempel:  
Om Du anger talet 3,4 och signifikansen 1 visas 3 som resultat.  
Om Du anger talet -6 och signifikansen -5 visas -10 som resultat.  
Om Du anger talet -0,6 och signifikansen -0,4 visas -0,8 som resultat.  
AVRUNDA.NEDÅT, AVRUNDA.UPPÅT, HELTAL, JÄMN, AVKORTA, RUNDA.UPP, AVRUNDA, UDDA  
TECKEN  
Med den här funktionen kan du beräkna ett tals förtecken (Sign).  
Funktionen returnerar 1 som resultat för ett positivt förtecken och -1 för ett negativt förtecken.  
Om talet är noll, ger funktionen också resultatet noll.  
Syntax:  
TECKEN( tal)  
tal är det tal vars förtecken Du ska bestämma.  
Exempel:  
Om Du anger talet 3,4 visas 1 som resultat.  
Om Du anger talet -4,5 visas -1 som resultat.  
ABS  
MAVRUNDA  
Resultatet är ett heltal som är den heltalsmultipel som ligger närmast talet av Multipel.  
Syntax  
MAVRUNDA( Tal;Multipel)  
Exempel  
Vilken heltalsmultipel av 3 ligger närmast talet 15,5?  
=MAVRUNDA( 15,5; 3) ger resultatet 15.  
ROT  
Om Du vill dra kvadratroten ur ett tal, anger Du talet i textfältet tal.  
Värdet för tal måste vara positivt.  
Syntax:  
ROT( tal)  
tal är det tal vars kvadratrot Du ska beräkna.  
Exempel:  
Kvadratroten för talet 16 är 4.  
Kvadratroten för talet -16 ger ett felmeddelande.  
ROT( ABS(-16)) = 4.  
UPPHÖJT.TILL, ABS  
ROTPI  
Resultatet är kvadratroten ur ett tal*PI.  
Syntax  
ROTPI( Tal)  
Exempel  
=ROTPI( 2) ger resultatet 2,506628.  
SLUMP.MELLAN  
Resultatet är ett slumptal som är ett heltal mellan Minsta tal och Största tal (båda inkluderade).  
För att beräkna på nytt trycker du på Skift+Ctrl+F9.  
Syntax  
SLUMP.MELLAN( Minsta tal;Största tal)  
Exempel  
=SLUMP.MELLAN( 20;30) ger ett heltal från 20 till 30 som resultat.  
SLUMP  
Med den här funktionen kan Du generera ett slumptal ur området 0 till 1.  
Dra upp ett område i tabellen, välj den här funktionen, markera fältet matris och klicka på OK.  
Det markerade området fylls med slumptal mellan 0 och 1.  
Syntax:  
SLUMP()  
ANTAL.OM  
Om Du vill räkna element som ska uppfylla vissa kriterier, anger Du det område som kriterierna ska tillämpas på i fältet område.  
Ange sökkriterierna i fältet kriterier.  
Syntax:  
ANTAL.OM( område; kriterier)  
område är det område som kriterierna ska tillämpas på.  
kriterier anger kriterierna i form av ett tal, ett uttryck eller en teckenföljd.  
Dessa kriterier bestämmer vilka celler som räknas.  
Ett sökkriterium kan t ex formuleras som 17, "17", ">100" eller "blå ".  
Du kan även skriva in en söktext som reguljärt uttryck, t ex "b.*" för alla ord som börjar på b.  
Du kan även ange ett cellområde som innehåller sökkriteriet.  
Exempel:  
Kriteriet 22,5 i området A1:E4 i exempeltabellen ska räknas.  
Ange A1:E4 i textfältet område och 22,5 som kriterium.  
1 visas som resultat.  
ANTAL.OM( A1:E4;22,5) ger 1.  
Ytterligare ett exempel finns vid SUMMA().  
ANTAL.TOMMA, SUMMA.OM.  
Kategorin Matris  
Här förklaras funktionerna inom kategorin Matris med hjälp av ett exempel.  
Till den här kategorin hör funktionerna ENHETSMATRIS, FREKVENS, MDETERM, MINVERT, MMULT, MTRANS, REGR, EXPREGR, PRODUKTSUMMA, SUMMAX2MY2, SUMMAX2PY2, SUMMAXMY2, TREND och EXPTREND.  
De beskrivs nedan.  
Vad är en matris?  
I tabellberäkning är en matris ett sammanhängande område med celler som innehåller värden.  
Ett kvadratiskt område med t.ex. 3 rader och 3 kolumner blir då en 3 x 3-matris:  
A  
B  
C  
1  
7  
31  
33  
2  
95  
17  
2  
3  
5  
10  
50  
Den minsta matrisen som kan finnas är en 1 x 2 - eller 2 x 1-matris bestående av två angränsande celler.  
Vad är en matrisformel?  
En formel, som utvärderar de enskilda värdena i ett cellområde, kallas matrisformel.  
Skillnaden jämfört med andra formler är att formeln inte bearbetar ett enskilt värde utan flera värden samtidigt.  
En matrisformel bearbetar inte bara flera värden utan kan även returnera flera värden.  
Resultatet av en matrisformel blir alltså i sin tur en matris.  
Det räcker med en enda matrisformel.  
Du väljer ett område med 3x3 celler på ett annat ställe, skriver in formeln "=10*A1:C3" och bekräftar med tangentkombinationen Kommando Ctrl +Skift+Retur.  
Resultat blir en 3 x 3-matris, där de enskilda värdena i cellområdet (A1:C3) multipliceras med 10.  
I %PRODUCTNAME Calc används operatorerna addition (+), subtraktion (-), multiplikation (*), division (/), exponent (^), kedjade tecken (&) och relationsoperatorer (=, <>, <, >, <=, >=).  
Operatorerna verkar på varje enskilt värde i cellområdet och returnerar resultatet i form av en matris om formeln angetts som en matrisformel.  
När jämförelseoperatorer används i matrisformler gäller samma regler för tomma celler som vid enkla jämförelser, d v s de tomma cellerna kan representera numeriskt 0 eller en tom sträng.  
Både matrisformeln {=A1:A2=""} och {=A1:A2=0} returnerar SANT om cellerna A1 och A2 är tomma.  
Matrisjämförelser med tomma celler beräknas på annat sätt i %PRODUCTNAME 5.0 än i tidigare versioner.  
När ska jag använda matrisformler?  
Om beräkningsförutsättningarna, d.v.s. formeln, ändras behöver du bara ändra på ett ställe.  
Då markerar du först hela matrisområdet och gör sedan den nödvändiga ändringen i matrisformeln.  
Matrisformler är dessutom ett utrymmesbesparande alternativ när flera värden ska utvärderas eftersom det inte behöver så mycket minne.  
I %PRODUCTNAME Calc finns det olika matematiska funktioner för beräkning med matriser, t.ex. funktionen MMULT som multiplicerar två matriser eller funktionen PRODUKTSUMMA som returnerar en skalärprodukt av två matriser.  
Matrisformler i %PRODUCTNAME Calc  
Du kan naturligtvis även skapa "normala" formler, där du anger områdesreferenser som parameterarna i en matrisformel.  
Resultatet bildas istället genom att referensområdet korsas med den rad eller kolumn, där formeln står.  
Om det inte finns någon korsning eller om området i korsningen omfattar flera kolumner eller rader returneras ett #Värde! som fel.  
I tidigare versioner av %PRODUCTNAME skapades en matris automatiskt när de ovannämnda operatorerna användes som parameter för en områdesreferens.  
Formeln "=Summa(B8 -(B10:B12))" returnerade automatiskt summan (B8-B10)+(B8-B11)+(B8-B12).  
Fr o m %PRODUCTNAME 5.0 gäller inte detta längre.  
En formel måste uttryckligen definieras som en matrisformel enligt mönstret {"=Summa(B8 -(B10:B12))"} för att det angivna cellområdet ska gälla som parameter.  
Om Du importerar tabelldokument som skapats i tidigare versioner av %PRODUCTNAME och där "normala" formler använts med cellområden som parametrar måste Du manuellt skapa matrisformler av de befintliga formlerna om Du vill få samma resultat.  
Då gör Du på följande sätt:  
Placera markören i den cell som innehåller den formel som ska konverteras och tryck på funktionstangenten F2.  
Tryck på Vänsterpil så flyttas markören ett steg åt vänster.  
Bekräfta formeln med kortkommandot Kommando Ctrl +Skift+Retur.  
Nu är formeln en matrisformel.  
Så här skapar du en matrisformel  
Om du skapar en matrisformel med Funktionsautopiloten måste du alltid markera rutan Matris om du vill få resultatet i form av en matris. (I annat fall returneras bara värdet i den vänstra övre cellen i den beräknade matrisen som resultat.)  
Om Du skriver in en matrisformel direkt i en cell så måste Du avsluta med Skift + Kommando Ctrl +Retur.  
Endast då gäller formeln som matrisformel.  
Matrisformler i %PRODUCTNAME Calc omges av klammerparentes.  
Du kan dock inte skapa en matrisformel genom att själv skriva in klammerparentestecknen eftersom %PRODUCTNAME Calc tolkar dem som text.  
Cellerna i en resultatmatris skyddas automatiskt mot ändringar.  
Men du kan ändra eller kopiera matrisformeln.  
Då måste du markera hela cellområdet, d.v.s. hela matrisen.  
Så här ändrar du en matrisformel  
Markera det cellområde eller den matris som innehåller matrisformeln.  
Tryck antingen på F2 eller placera markören på inmatningsraden.  
Båda alternativen har samma effekt.  
Nu kan du redigera formeln.  
När du har gjort ändringar bekräftar du med kortkommandot Kommando Ctrl +Skift+Retur.  
Du kan formatera de enskilda delarna i en matris på olika sätt (t.ex. ge dem olika teckensnittsfärger).  
Du behöver bara markera det önskade cellområdet och tilldela det önskade attribut.  
Så här kopierar du en matrisformel  
Markera det cellområde eller den matris som innehåller matrisformeln.  
Tryck på F2 eller placera markören på inmatningsraden.  
Kopiera formeln från inmatningsraden med Kommandot Ctrl +C.  
Markera det cellområde där matrisformeln ska infogas, och tryck åter på F2 eller placera markören på inmatningsraden.  
Klistra in formeln från urklippet på inmatningsraden med Kommando Ctrl +V och bekräfta med Kommando Ctrl +Skift+Retur.  
Nu får det nya markerade området en matrisformel.  
Så här anpassar du ett matrisområde  
Om Du vill ändra storleken på en resultatmatris, t ex om matrisformeln innehåller ett område som Du vill dölja, gör Du på följande sätt:  
Markera det cellområde eller den matris som innehåller matrisformeln.  
Till höger nedtill i det markerade området finns en liten markering, som Du kan dra i med musen om Du vill förstora eller förminska området.  
Observera att själva matrisformeln inte ändras när Du anpassar matrisområdet.  
Anpassningen påverkar bara det område där resultatet visas.  
Om Du håller Ctrl nedtryckt när Du drar så skapas en kopia av matrisformeln i det markerade området.  
ENHETSMATRIS  
Bestämmer den kvadratiska enhetsmatrisen för en bestämd storlek.  
Enhetsmatrisen är en kvadratisk matris, där huvuddiagonalelementen är lika med 1 och alla andra matriselement är lika med 0.  
Syntax  
ENHETSMATRIS( dimension)  
dimension bestämmer storleken för enhetsmatrisen.  
Exempel  
Markera ett kvadratiskt område i tabellen, t ex från A1 till E5.  
Öppna funktionen ENHETSMATRIS utan att upphäva markeringen.  
Markera rutan Matris.  
Ange dimensionen för den önskade enhetsmatrisen, i det här fallet 5.  
Klicka på OK.  
Du kan även skriva in formeln =Enhetsmatris (5) i den sista cellen i det markerade området (i det här fallet E5) och avsluta kommandot med Skift+Kommando+Retur Skift+Ctrl+Retur.  
Nu visas enhetsmatrisen i området A1:E5.  
FREKVENS  
Returnerar en frekvensfördelning som en matris i en kolumn.  
Inom en given mängd värden och ett givet antal intervaller eller klasser beräknas vilket antal värden som ligger inom de enskilda intervallerna.  
Syntax  
FREKVENS( data; klasser)  
data är en matris eller referens till den mängd värden som ska beräknas.  
klasser är en matris för klassindelning.  
Exempel  
Observera följande data.  
I kolumn A står mätvärden (data) i valfri ordningsföljd.  
I kolumn B har Du angett de övre gränserna för de klasser som Du vill dela in data i.  
Värdet 5 i cell B1 innebär att Du vill att det första resultatet av funktionen FREKVENS ska ange det antal mätvärden (data) som är mindre än eller lika med 5.  
I B2 står talet 10 som nästa klassgräns.  
Det andra resultatet av funktionen FREKVENS ska alltså ange det antal mätvärden som är större än 5 och mindre än eller lika med 10.  
I cell B6 har Du skrivit in texten ">25" som orientering.  
A  
B  
C  
1  
12  
5  
1  
2  
8  
10  
3  
3  
24  
15  
2  
4  
11  
20  
3  
5  
5  
25  
1  
6  
20  
>25  
1  
7  
16  
8  
9  
9  
7  
10  
16  
11  
33  
Markera ett område i en kolumn där frekvenserna ska anges (Du måste markera ett fält mer än det finns övre klassgränser för de värden som ligger över den sista klassgränsen).  
I det här exemplet markerar du området C1:C6.  
Öppna funktionen FREKVENS i Funktionsautopiloten.  
Välj sedan en kolumn, där du skrivit in klassgränserna (B1:B6), som klasser.  
Markera Matris och klicka på OK.  
Nu visas frekvensberäkningen i det ursprungligen markerade området C1:C6.  
ANTAL, DANTAL.  
MDETERM  
Returnerar determinanten för en kvadratisk matris.  
Du behöver inte definiera något utdataområde.  
Syntax  
MDETERM( matris)  
matris är den kvadratiska matris, vars determinant ska bestämmas.  
Exempel  
MDETERM( C3:D4) = -6.  
MINVERT, MMULT, MTRANS.  
MINVERT  
Beräknar inversen för en matris (omvänd matris).  
Den inverterade matrisen är den matris som, multiplicerad med ursprungsmatrisen, ger enhetsmatrisen.  
Syntax  
MINVERT( matris)  
matris är den kvadratiska matris, som ska inverteras.  
Exempel  
Markera ett kvadratiskt område och öppna den här funktionen.  
Markera utgångsmatrisen, markera rutan Matris och klicka på OK.  
INDEX, MMULT.  
MMULT  
Beräknar produkten av två matriser.  
Den kvadratiska resultatmatrisen har samma antal rader och kolumner.  
Syntax  
MMULT( matris 1; matris 2)  
matris 1 är den första matrisen för matrisprodukten.  
matris 2 är den andra matrisen med samma antal rader.  
Exempel  
Markera t.ex. ett kvadratiskt område.  
Öppna den här funktionen.  
Välj först den ena matrisen 1 och sedan den andra matrisen 2.  
Markera rutan Matris i Funktionsautopiloten.  
Klicka på OK.  
Resultatmatrisen visas i det område som du markerade först.  
MDETERM, MINVERT, MTRANS.  
MTRANS  
Här kan Du byta ut (transponera) rader och kolumner i en matris.  
Syntax  
MTRANS( matris)  
matris är den matris i en tabell som ska transponeras.  
Exempel  
Markera ett område som kan rymma den transponerade matrisen.  
Om ursprungsmatrisen består av n antal rader och m antal spalter måste det markerade området innehålla minst m antal rader och n antal spalter.  
Skriv in formeln direkt, välj ursprungsmatrisen och tryck på Skift+Kommando+Retur Skift+Ctrl+Retur.  
Om du använder Funktionsautopiloten markerar du rutan Matris.  
Den transponerade matrisen visas i det markerade målområdet.  
Cellerna i den transponerade matrisen skyddas automatiskt mot ändringar.  
MDETERM, MINVERT, MMULT.  
REGR  
Beräknar en linje som visar den bästa linjära regressionsanpassningen för givna data och ger som resultat en matris, vars element beskriver linjen.  
Syntax  
REGR( data_y; data_x; typ_av_linje; statistik)  
data_y är matrisen med y-data.  
data_x (valfri) är matrisen med x-data.  
typ_av_linje (valfri).  
Om linjen ska gå genom nollpunkten, anger du linjetyp = 0.  
statistik (valfri).  
Om statistik = 0 så beräknas bara regressionskoefficienterna.  
Annars visas ytterligare statistikvärden.  
Exempel  
Den här funktionen returnerar en matris. (Den ska alltså behandlas som övriga matrisfunktioner enligt beskrivningen i sidans inledning.) Markera det område där svaren ska visas.  
Öppna den här funktionen.  
Välj y-data.  
Ange fler parametrar om du vill.  
Markera Matris och klicka på OK.  
Som resultat visas minst (om statistik = 0) lutningen för regressionslinjen och skärningspunkten mot Y-axeln.  
Om statistik inte är lika med noll visas fler resultat.  
Ytterligare resultat för REGR-funktionen:  
Titta på följande exempel:  
A  
B  
C  
D  
E  
F  
G  
1  
x1  
x2  
y  
REGR-värden  
2  
4  
7  
100  
4,17  
-3,48  
82,33  
3  
5  
9  
105  
5,46  
10,96  
9,35  
4  
6  
11  
104  
0,87  
5,06  
#Saknas  
5  
7  
12  
108  
13,21  
4  
#Saknas  
6  
8  
15  
111  
675,45  
102,26  
#Saknas  
7  
9  
17  
120  
8  
10  
19  
133  
I kolumn A visas några X1-värden, i kolumn B visas några X2-värden och i kolumn C visas Y-värdena.  
Alla de här värdena har du redan lagt in i tabellen.  
Funktionen REGR kräver att du kryssar för rutan Matris i Funktionsautopiloten.  
På sidan 2 i Funktionsautopiloten väljer du nu följande värden i tabellen (eller matar in dem via tangentbordet):  
data_y är C2:C8  
data_x är A2:B8  
typ_av_linje och statistik har båda satts till lika med 1.  
När du klickar på OK fyller %PRODUCTNAME Calc i de synliga REGR-värdena i exemplet ovan.  
För varje cell i REGR-matrisen är formeln i formellisten {=REGR(C2:C8;A2:B8;1;1)}.  
De beräknade REGR-värdena betyder följande:  
E2 och F2:  
Lutningen m för regressionslinjen y=b+m*x för värdena x1 och x2.  
Värdena returneras i omvänd ordning, d.v.s. lutningen för x2 i E2 och lutningen för x1 i F2.  
G2:  
Skärningspunkten b mot Y-axeln.  
E3 och F3:  
Standardskattningsfel för lutningsvärdena.  
G3:  
Standardskattningsfel för axelavsnittet.  
E4:  
Korrelationskoefficienten.  
F4:  
Standardskattningsfel för Y-värdena som beräknats från regressionen.  
E5:  
F-värdet från variansanalysen.  
F5:  
Frihetsgraderna från variansanalysen.  
E6:  
Summan av de kvadratiska avvikelserna för de skattade y-värdena från det aritmetiska medelvärdet.  
F6:  
Summan av de kvadratiska avvikelserna för de skattade y-värdena från de givna y-värdena.  
EXPREGR, TREND, EXPTREND.  
EXPREGR  
Den här funktionen beräknar en exponentialkurva som passar givna data (exponentiell regression, y=b*m^x).  
Syntax  
EXPREGR( data_y; data_x; typ_av_funktion; statistik)  
data_y är matrisen med y-data.  
data_x (valfri) är matrisen med x-data.  
typ_av_funktion (valfri).  
I annat fall beräknas även funktionerna y = b*m^x.  
statistik (valfri).  
Om statistik = 0 så beräknas bara regressionskoefficienterna.  
Exempel  
Se REGR.  
Inga kvadratsummor returneras som resultat.  
REGR, TREND, EXPTREND.  
PRODUKTSUMMA  
Summerar produkterna av argument i matriser.  
Detta innebär alltså en summa av produkter.  
Syntax  
PRODUKTSUMMA( matris 1; matris 2...matris 30)  
matris 1, matris 2...matris 30 är matriser, vars argument ska multipliceras.  
Exempel  
=PRODUKTSUMMA( C3;D6;D8;D3) ger resultatet 270.  
MMULT, PRODUKT, SUMMA.  
SUMMAX2MY2  
Summerar skillnaden mellan kvadraterna för motsvarande värden i två matriser.  
Detta innebär alltså en summa av skillnaderna mellan kvadraterna.  
Syntax  
SUMMAX2MY2( matris _x; matris_y)  
matris_x är den första matrisen, vars element ska kvadreras och adderas.  
matris_y är den andra matrisen, vars element ska kvadreras och subtraheras.  
Exempel  
=SUMMAX2MY2( D6; D8) ger resultatet -27.  
PRODUKTSUMMA, SUMMAX2PY2, SUMMAXMY2.  
SUMMAX2PY2  
Summan av kvadraterna i två matriser adderas.  
Syntax  
SUMMAX2PY2( matris_x; matris_y)  
matris_x är den första matrisen, vars argument ska kvadreras och summeras.  
matris_y är den andra matrisen, vars argument ska kvadreras och summeras.  
Exempel  
=SUMMAX2PY2( D6;D8) ger resultatet 45.  
PRODUKTSUMMA, SUMMAX2MY2, SUMMAXMY2.  
SUMMAXMY2  
Summerar kvadraterna på skillnaden mellan två matriser.  
Syntax  
SUMMAX2MY2( matris_x; matris_y)  
matris_x är den första matrisen, vars element ska subtraheras och kvadreras.  
matris_y är den andra matrisen, vars element ska subtraheras och kvadreras.  
Exempel  
=SUMMAXMY2( C4;C9) ger resultatet 64.  
PRODUKTSUMMA, SUMMAX2MY2, SUMMAX2PY2.  
TREND  
Beräknar värden som erhålls längs en linjär trend.  
Syntax  
TREND( data_y; data_x; nya_data_x; typ_av_linje)  
data_y är matrisen med y-data.  
data_x (valfri) är matrisen med x-data.  
nya_data_x (valfri) är matrisen med X-data som används för ny beräkning av värden.  
typ_av_linje (valfri).  
I annat fall beräknas även förskjutna linjer.  
Standardinställningen för typ är <> 0.  
Exempel  
Markera ett område där trenddata ska visas.  
Öppna den här funktionen.  
Ange området med utgångsdata eller markera det med musen.  
Markera rutan Matris.  
Klicka på OK.  
Nu visas de trenddata som beräknats från utgångsdata.  
REGR, EXPREGR, EXPTREND.  
EXPTREND  
Beräknar punkter på en exponentiell regressionsfunktion i en matris.  
Syntax  
EXPTREND( data_y; data_x; nya_data_x; typ_av_funktion)  
data_y är matrisen med y-data.  
data_x (valfri) är matrisen med x-data.  
nya_data_x (valfri) är matrisen med x-data som används för ny beräkning av värden.  
typ_av_funktion (valfri).  
I annat fall beräknas även funktionerna y = b*m^x.  
Exempel  
Den här funktionen returnerar en matris. (Den ska alltså behandlas som de andra matrisfunktionerna enligt beskrivningen i sidans inledning.) Markera ett område där svaren ska visas.  
Öppna den här funktionen.  
Välj Y-data.  
Ange fler parametrar om du vill.  
Markera Matris och klicka på OK.  
REGR, EXPREGR, TREND.  
Kategorin Statistik  
Här visas med ett exempel de funktioner som står till förfogande i kategorin Statistik.  
Det rör sig om följande funktioner:  
SKÄRNINGSPUNKT, ANTAL, ANTALV, B, RKV, BETAINV, BETAFÖRD, BINOMFÖRD, CHI2INV, CHI2TEST, CHI2FÖRD, EXPONFÖRD,  
FINV, FISHER, FISHERINV, FTEST, FFÖRD, GAMMAINV, GAMMALN, GAMMAFÖRD, GAUSS, GEOMEAN, TRIMMEDEL, ZTEST, HARMMEDEL, HYPGEOMFÖRD,  
STÖRSTA, MINSTA, KONFIDENS, KORREL, KOVAR, KRITBINOM, TOPPIGHET, LOGINV, LOGNORMFÖRD,  
MAX, MAXA, MEDIAN, MIN, MINA, MEDELAVV, MEDEL, MEDELA, TYPVÄRDE, NEGBINOMFÖRD, NORMINV, NORMFÖRD, PEARSON, PHI, POISSON, PERCENTIL, PROCENTRANG, KVARTIL,  
RANG, SNEDHET, PREDIKTION, STDAV, STDAVA, STDAVP, STDAVPA, STANDARDISERA, NORMSINV, NORMSFÖRD, LUTNING, STDFELYX, KVADAVV, TINV, TTEST, TFÖRD, VARIANS, VARIANSA, VARIANSP, VARIANSPA, PERMUT, PERMUT2, SANNOLIKHET, WEIBULL.  
Funktionerna beskrivs i följande underkapitel.  
Statistikfunktioner i analys-add-in  
Några exempel går bara att förklara med hjälp av en tabell.  
Använd i sådana fall följande tabell som utgångspunkt.  
C  
D  
2  
x-värde  
y-värde  
3  
-5  
-3  
4  
-2  
0  
5  
-1  
1  
6  
0  
3  
7  
2  
4  
8  
4  
6  
9  
6  
8  
De omfattande statistikfunktionerna beskrivs i följande underkapitel:  
Kategorin Tabell  
Här visas med ett exempel de funktioner som står till förfogande i kategorin Tabell.  
Det rör sig om följande funktioner:  
ADRESS, OMRÅDEN, DDE, FELTYP, INDEX, INDIREKT, KOLUMN, KOLUMNER, LETARAD, TABELL, TABELLER, PASSA;, FÖRSKJUTA, LETAUPP, FORMATMALL, VÄLJ, LETAKOLUMN, RAD och RADER.  
De beskrivs nedan.  
ADRESS  
Anger en cells adress (referensen) om Du anger radnumret och kolumnnumret.  
Som ett alternativ kan Du bestämma om adressen ska visas absolut (t ex i formen $A$1) eller relativt (som A1) eller blandat (A$1 eller $A1).  
Du kan också ange tabellens namn.  
Syntax  
ADRESS( rad; kolumn; ABS; tabell)  
rad är cellreferensens radnummer.  
kolumn är cellreferensen kolumnnummer (inte bokstaven)  
ABS bestämmer typen av referens:  
1 eller tom:  
Absolut ($A$1)  
2:  
Rad absolut, kolumn relativ (A$1)  
3:  
Rad relativ, kolumn absolut ($A1)  
4:  
Relativ (A1)  
tabell är namnet på en tabell.  
Exempel  
Tabell2.A$1  
Sätt t.ex. den här funktionen i cellen B2.  
Om värdet -6 står i tabell2.  
A1, kan du via funktionen i B2 indirekt hänvisa till cellen som det refererats till på detta sätt, genom att t.ex. skriva =ABS( INDIREKT(B2)) i en formel.  
Du får därmed cellinnehållets absolutbelopp för cellen vars adress har angetts i B2, i detta fall 6.  
KOLUMN, RAD.  
OMRÅDEN  
Anger antalet områden som tagits upp inom en referens.  
Ett område (delområde) kan bestå av flera sammanhängande celler (cellområde) eller av en enda cell.  
Syntax  
OMRÅDEN( referens)  
referens är en referens till en cell eller ett cellområde.  
Exempel  
=OMRÅDEN( A1:B3;F2;G1) returnerar 3 eftersom tre områden räknas upp här.  
=OMRÅDEN( Alla) returnerar 1, om du har definierat ett område med namnet Alla innan dess i Data - Definiera område.  
Referenser till raderade områden (t.ex. refererade tabeller eller kolumner) importeras och exporteras av %PRODUCTNAME.  
ADRESS, INDEX, KOLUMN, KOLUMNER, RAD, RADER.  
DDE  
Returnerar resultatet för en DDE-operator.  
Om innehållet i det länkade området ändras, ändras också det värde som formeln returnerar.  
Syntax  
DDE( server;fil;område;läge)  
server är namnet på ett serverprogram. %PRODUCTNAME -programmen har servernamnet "Soffice":  
fil är namnet på filen, inklusive dess fullständiga sökväg.  
område är ett område ur vilket data ska läsas.  
Läge är en valfri parameter som styr hur data omvandlas till tal av DDE-servern. (Denna parameter är ny.  
Ifall Du vill öppna tabellen med en föregående version av %PRODUCTNAME Calc, bör Du avstå från denna parameter.)  
Läge  
Effekt  
0 eller saknas  
Talformat ur "standard "-cellformatmallen  
1  
Data tolkas alltid med standardformatet för engelska (US)  
2  
Data övertas som text, ingen omvandling till tal  
Exempel  
=DDE( "soffice" ;"c:\office5\document\data1.sdc" ;"Tabelle1.A1") läser innehållet i cellen A1 i tabell 1 i %PRODUCTNAME Calc-dokumentet Data1.sdc.  
=DDE( "soffice" ;"c:\office5\document\Motto.sdw" ;"Dagensmotto") ger dagens motto som innehåll i den cell i vilken denna formel står.  
Förutsättningen är att Du har skrivit in det på en rad i %PRODUCTNAME Writer-dokumentet Motto.sdw, och att denna rad är den första raden i det namngivna området (%PRODUCTNAME Writer-menyn Infoga-Område...) Så snart dagens motto ändras i %PRODUCTNAME Writer-dokumentet och sparas på nytt, är det tillgängligt i alla de %PRODUCTNAME Calc-celler i vilka denna DDE-länk har definierats.  
FELTYP  
Denna funktion returnerar numret på en felkod som uppträtt i en annan cell i form av ett värde.  
Med hjälp av detta nummer kan Du visa en egen feltext.  
Den fördefinierade felkoden från %PRODUCTNAME Calc visas i statuslisten när Du klickar på cellen med felet.  
Syntax  
FELTYP( referens)  
referens är en referens till en cell i vilken ett fel har rapporterats.  
Exempel  
Om det t ex står Err:518 i cellen A1, ger funktionen =FELTYP( A1) värdet 518.  
ÄRREF, ÄRF, ÄRFEL, ÄRFORMEL.  
ÄREJTEXT, ÄRTOM, ÄRLOGISK, ÄRSAKNAD, ÄRTEXT, ÄRTAL.  
INDEX  
INDEX ger innehållet i en cell, som har definierats med radnummer och kolumnnummer och i förekommande fall av området.  
Syntax  
INDEX( referens;rad;kolumn;område)  
referens är en referens till celler via direkt skrivsätt eller genom att namnet på ett område har angetts.  
Om referensen är ett multipelområde ska den stå inom runda parenteser, även när Du nämner den med namn.  
rad (valfri) är numret på den rad i det område som nämns i referensen.  
kolumn (valfri) är numret på den kolumn i det område som nämns i referensen.  
område (valfri) är en parameter som betecknar delområdets index om det finns mer än ett område inom det område som det refererats till.  
Exempel  
=INDEX( Priser;4;1) ger värdet som står på rad 4 och kolumn 1 i databasområdet som du har försett med namnet Priser under Data - Definiera område.  
=INDEX( Summor;4;1) ger värdet som står på rad 4 och kolumn 1 i området med namnet Summor som du har tilldelat under Infoga - Namn - Definiera....  
=INDEX( Multipel;4;1) ger värdet som står på rad 4 och kolumn 1 i multipelområdet som du har försett med namnet Multipel under Infoga - Namn - Definiera....  
Multipelområdet kan bestå av flera rektangulära cellområden, som vart och ett kan ha en rad 4 och en kolumn 1.  
Om du vill anropa det andra blocket i detta multipelområde anger du 2 som sista parameter område.  
=INDEX( A1:B6;1,1) anger värdet uppe till vänster i området A1:B6.  
LETARAD, PASSA, LETAUPP, VÄLJ, LETAKOLUMN.  
INDIREKT  
Ger tillbaka den referens som står i den cell eller det cellområde som Du har angett med argumentet referens.  
Den här funktionen kan också skapa ett område ur en motsvarande teckenföljd.  
Syntax  
INDIREKT( referens)  
referens är den cell eller det område vars innehåll ska utvärderas. referens ges i textformat.  
Exempel  
=INDIREKT( A1) ger 100, när referensen C108 står i A1 och värdet 100 står i cell C108.  
=SUMMA( INDIREKT("a1: "& ADRESS(1;3))) summerar cellerna i området från A1 till den cell vars adress är definierad genom rad 1 och kolumn 3.  
Det är alltså området A1:C1 som summeras.  
FÖRSKJUTA.  
KOLUMN  
Returnerar kolumnnumren för en referens.  
Ifall ett cellområde är parameter, sker utmatningen av de tillhörande kolumnnumren i en enradig matris om formeln skrivs in som en matrisformel.  
Om funktionen KOLUMN med en områdesreferens som parameter inte används i en matrisformel, så fastställs endast kolumnnumret för områdets första cell.  
Syntax  
KOLUMN( referens)  
referens är referensen till ett cellområde vars kolumnnummer ska räknas fram.  
Argumentet kan också vara en enstaka cell.  
Om Du inte anger någon referens, så fastställs kolumnnumret för den cell i vilken formeln matas in. %PRODUCTNAME Calc sätter automatiskt referensen till den aktuella cellen.  
Exempel  
=KOLUMN( B3) ger 2, eftersom kolumn B är den andra kolumnen i tabellen.  
{=KOLUMN(D3:G10)} ger den enradiga matrisen (4, 5, 6, 7), eftersom kolumnerna D till G är den fjärde till sjunde kolumnen i tabellen.  
=KOLUMN( D3:G10) ger 4 eftersom kolumn D är tabellens fjärde kolumn och funktionen KOLUMN inte används som matrisformel. (I detta fall tas alltid matrisens första värde som resultat.)  
{=KOLUMN(B2:B7)} och =KOLUMN(B2:B7) ger båda 2 eftersom referensen bara innehåller kolumn B som tabellens andra kolumn. (Eftersom det hos enspaltiga områden bara finns ett kolumnnummer, gör det här inte någon skillnad om formeln används som matrisformel eller inte.)  
=KOLUMN() ger 3 om formeln har matats in i kolumn C.  
{=KOLUMN(hare)} ger den enradiga matrisen (3, 4) om "hare "är det namngivna området (C1:D3).  
Funktionen KOLUMN är inte kompatibel med tidigare %PRODUCTNAME -versioner.  
När Du laddar äldre %PRODUCTNAME Calc-dokument, bör Du tänka på att KOLUMN() hittills har returnerat resultaten i en lodrät enspaltig m x 1-matris i stället för i en vågrät enradig 1 x n-matris.  
KOLUMNER, RAD.  
KOLUMNER  
Returnerar antalet kolumner i en referens.  
Syntax  
KOLUMNER( matris)  
matris är referensen till ett cellområde vars kolumnantal ska uträknas.  
Argumentet kan också vara en enda cell.  
Exempel  
=Kolumner( B5) ger 1 eftersom en cell bara omfattar en kolumn.  
=KOLUMNER( A1:C5) returnerar 3, eftersom referensen omfattar tre kolumner.  
=KOLUMNER( hare) ger 2 om "hare "är det namngivna området (C1:D3).  
Funktionen KOLUMNER visar fr o m %PRODUCTNAME 5.0 ett annat tolkningssätt än i tidigare versioner om Du överlämnar en internt genererad matris som parameter.  
När Du laddar äldre %PRODUCTNAME Calc-dokument och har använt sådana parametrar, bör Du tänka på att KOLUMNER() i sådana fall nu returnerar andra resultat (inte radernas antal som tidigare, utan kolumnernas).  
KOLUMN, RADER.  
LETARAD  
Lodrät sökning och hänvisning till höger därom liggande celler.  
Funktionen returnerar då värdet för en viss kolumn i matrisen på samma rad som namngetts med index.  
Syntax  
=LETARAD( sökkriterium;matris;index;sorterad)  
sökkriterium är värdet som ska sökas i matrisens första kolumn.  
matris är referensen som ska bestå av minst två kolumner.  
index är numret på den kolumn inom matrisen i vilken det returnerade värdet står.  
Den första kolumnen har nummer 1.  
sorterad är en valfri parameter, som anger om den första kolumnen i matrisen är sorterad i stigande ordning (detta är standard).  
Ange här det logiska värdet FALSK om den första kolumnen inte är sorterad i stigande ordning.  
Det går mycket snabbare att söka igenom sorterade kolumner, och funktionen returnerar alltid ett värde, även om det exakta sökvärdet inte har hittats (såvida det ligger mellan det största och minsta värdet i den sorterade listan).  
I osorterade listor måste det exakta sökvärdet hittas, annars returnerar funktionen felet värde ej tillgängligt.  
Exempel  
Du vill mata in numret på en rätt på matsedeln (i cell A1), varefter namnet på rätten omedelbart ska visas i form av text i cellen bredvid (B1).  
Tilldelningen av nummer till namn står i matrisen D1:E100.  
I D1 står t.ex. 100 och i E1 står namnet Grönsakssoppa osv för 100 rätter.  
Du behöver alltså inte använda den valfria parametern sorterad.  
Infoga följande formel i B1:  
=LETARAD( A1; D1:E100; 2)  
Så snart Du skriver in ett nummer i A1 visas den därtill hörande texten i B1, vilken står i den andra kolumnen till referensen D1:E100.  
Om Du skriver in ett icke-existerande nummer visas texten med det närmast lägre numret.  
Då visas ett felmeddelande om ett icke-existerande nummer skrivs in.  
INDEX, PASSA, LETAUPP, LETAKOLUMN.  
Tabell  
Bestämmer tabellnumret för en referens eller en teckensträng som är ett tabellnamn.  
Om Du inte har angett någon parameter, så returneras tabellnumret för den tabell i vilken formeln står.  
Syntax  
Tabell( referens)  
referens är valfri och är referensen till en cell, ett område eller ett tabellnamns teckensträng.  
Exempel  
=TABELL( Tabell2.A1) ger 2 om Tabell2 är andra tabellen i ordningsföljden.  
Tabeller  
Bestämmer antalet tabeller för en referens.  
Om ingen parameter är angiven, returneras antalet tabeller i det aktuella dokumentet.  
Syntax  
Tabeller( referens)  
referens är referensen till en cell eller ett område.  
Denna parameter är valfri.  
Exempel  
=TABELLER( Tabell1.A1:Tabell3.G12) ger 3 om tabellerna Tabell1, Tabell2 och Tabell3 existerar i denna ordningsföljd.  
PASSA  
Bestämmer en position i en matris efter en värdejämförelse.  
Funktionen returnerar det påträffade värdets position i sökmatrisen i form av ett tal.  
PASSA( sökkriterium;sökmatris;typ)  
sökkriterium är det värde som Du vill söka efter i enrads - eller enkolumnsmatrisen.  
sökmatris är den referens i vilken sökningen utförs.  
typ kan anta värdena 1, 0 eller -1.  
Vid typ = -1 antas att sorteringen är fallande. (Funktionen har ändrats i %PRODUCTNAME 6.0 och motsvarar nu funktionen med samma namn i Microsoft Excel.)  
Om typ = 0 måste en exakt överensstämmelse hittas.  
Om sökkriteriet hittas flera gånger returnerar funktionen den första sökträffen.  
Bara vid typ = 0 är en sökning med reguljära uttryck tillåten.  
Om typ = 1 eller om den tredje parametern saknas, returneras det sista värdet som är mindre eller lika med sökkriteriet.  
Detta gäller även om sökmatrisen inte är sorterad.  
För typ = -1 returneras det första värdet som är större eller lika med sökkriteriet.  
Exempel  
=PASSA( 200; D1:D100) söker igenom området D1:D100, som sorterats enligt kolumn D, efter förekomster av värdet 200.  
Så snart detta värde har påträffats returneras radnumret för den rad där värdet hittats.  
Om ett högre värde påträffades vid sökningen i kolumnen, returneras numret på den föregående raden.  
INDEX, LETARAD, LETAKOLUMN.  
FÖRSKJUTA  
Returnerar värdet för en cell som är förskjuten ett visst antal rader och kolumner jämfört med en annan cell.  
Syntax  
FÖRSKJUTA( referens;rader;kolumner;höjd;bredd)  
referens är den cell från och med vilken funktionen beräknar den nya referensen.  
rader är det antal rader med vilken referensen förskjuts uppåt (negativt värde) eller nedåt.  
kolumner är antalet rader med vilket referensen förskjuts åt vänster (negativt värde) eller höger.  
höjd är den vertikala höjden, som Du kan ange om Du vill, för ett område som börjar vid den nya referenspositionen.  
bredd är den horisontella bredden, som Du kan ange om Du vill, för ett område som börjar vid den nya referenspositionen.  
Exempel  
=FÖRSKJUTA( A1; 2, 2) returnerar värdet i cell C3 (A1 förskjuten med två rader och två kolumner snett nedåt åt höger).  
Om 100 står i C3 ger denna funktion värdet 100 som resultat.  
=SUMMA( FÖRSKJUTA(A1; 2; 2; 5; 6)) bestämmer summan av området som börjar vid cell C3 och som är 5 rader högt och 6 kolumner brett, d.v.s. området C3:H7.  
LETAUPP  
Funktionen returnerar innehållet i en cell, som letas upp på en rad eller i en kolumn med ett sökkriterium.  
Om Du vill kan Du låta det tilldelade värdet (med samma index) returneras till en annan rad eller en annan kolumn.  
De behöver inte ligga bredvid varandra.  
För LETAUPP gäller det dessutom att sökvektorn måste vara sorterad, eftersom sökningen annars inte ger några användbara resultat.  
Syntax  
LETAUPP( sökkriterium;sökvektor;resultatvektor)  
sökkriterium är det värde som sökningen gäller, och vilket Du har angett direkt eller som referens.  
sökvektor är det enradiga eller enspaltiga område i vilket sökningen ska utföras.  
resultatvektor är ett annat enradigt eller enspaltigt område ur vilket funktionens resultat hämtas.  
Resultatet är den cell i resultatvektorn som har samma index som fyndplatsen i sökvektorn.  
Exempel  
=LETAUPP( A1; D1:D100;F1:F100) letar upp den cell i området D1:D100 som motsvarar det tal som Du anger i A1.  
Indexet till fyndplatsen tas fram, om det t ex är den 12:e cellen i området.  
Därefter returneras innehållet i den 12:e cellen i resultatvektorn som ett funktionsvärde.  
INDEX, LETARAD, LETAKOLUMN.  
FORMATMALL  
Tilldelar formelcellen en formatmall.  
Efter ett inställbart tidsintervall kan en annan formatmall tilldelas.  
På så sätt kan du med addition lägga till funktionen till en annan funktion, utan att ändra dess värde.  
Exempel: =.. .+FORMATMALL( OM(AKTUELL()>3 ;"röd" ;"grön")) färgar cellen med mallen "röd "om värdet är större än 3.  
Båda cellformaten "röd" och "grön "måste vara definierade innan.  
Syntax  
FORMATMALL( formatmall;tid;formatmall2)  
formatmall1 är namnet på en cellformatmall som tilldelas cellen.  
Namnen på mallarna ska stå inom citattecken.  
tid är ett tidsintervall i sekunder, som Du kan ange om Du vill.  
Om den här parametern saknas byts formatmallen inte ut efter en viss tid.  
formatmall2 är namnet på en cellformatmall, som Du kan ange om Du vill, och som tilldelas cellen efter det att tidsintervallet har gått ut.  
Om denna parameter saknas sätts "Standard".  
Exempel  
Därefter får den formatet Standard.  
Båda cellformaten måste vara definierade innan.  
VÄLJ  
Returnerar det värde som bestämts ur ett index och som hämtats ur en lista på upp till 30 värden.  
Syntax  
VÄLJ( index;värde 1;...värde 30)  
Anger vilket värde som ska tas ur listan.  
Värde 1...Värde 30 är listan över de värden som har angetts som referens till en cell eller som ett eget värde.  
Exempel  
För A1 = 4 returnerar funktionen texten Idag.  
För A1 = 7 returnerar den innehållet i den första cellen i det namngivna området Idag.  
INDEX.  
Vågrät sökning och hänvisning till celler som ligger direkt nedanför.  
Den här funktionen kontrollerar om det står ett visst värde på den första raden i en matris.  
Funktionen returnerar då värdet för en viss rad i matrisen på samma rad som namngetts med index.  
Syntax  
=LETAKOLUMN( sökkriterium;matris;index;sorterad)  
Endast rader byts ut mot kolumner.  
INDEX, LETARAD, PASSA, LETAUPP.  
RAD  
Returnerar radnumren för en referens.  
Ifall ett cellområde är parameter, sker utmatningen av de tillhörande radnumren i en enspaltig matris om formeln skrivs in som en matrisformel.  
Om funktionen RAD med en områdesreferens som parameter inte används i en matrisformel, så fastställs endast radnumret för områdets första cell.  
Syntax  
RAD( referens)  
referens är referensen till ett cellområde vars radnummer ska fastställas.  
Argumentet kan också vara en enstaka cell.  
Ifall Du inte anger någon referens, så fastställs radnumret för den cell i vilken formeln matas in. %PRODUCTNAME Calc sätter automatiskt referensen till den aktuella cellen.  
Exempel  
=RAD( B3) ger 3 eftersom referensen hänvisar till tabellens tredje rad.  
{=RAD(D5:D8)} ger den enspaltiga matrisen (5, 6, 7, 8) eftersom den angivna referensen innehåller raderna 5 till 8.  
=RAD( D5:D8) ger 5 eftersom funktionen RAD inte används som matrisformel och därför returneras bara numret för referensens första rad.  
{=RAD(A1:E1)} och =RAD(A1:E1) ger båda 1 eftersom referensen bara innehåller rad 1 som tabellens första rad. (Eftersom det bara finns ett radnummer hos enradiga områden, gör det här inte någon skillnad om formeln används som matrisformel eller inte.)  
=RAD() ger 3 om formeln har matats in på rad 3.  
{=RAD(hare)} ger den enspaltiga matrisen (1, 2, 3) om "hare "är det namngivna området (C1:D3).  
Funktionen RAD är inte kompatibel med tidigare %PRODUCTNAME -versioner.  
När Du laddar äldre %PRODUCTNAME Calc-dokument, bör Du tänka på att RAD() hittills har returnerat resultaten i en vågrät enradig 1 x n-matris i stället för i en lodrät enspaltig m x 1-matris.  
KOLUMN, RADER.  
RADER  
Returnerar antalet rader i en referens.  
Syntax  
RADER( matris)  
matris är referensen till ett cellområde vars radantal ska fastställas.  
Argumentet kan också vara en enda cell.  
Exempel  
=Rader( B5) ger 1 eftersom en cell bara omfattar en rad.  
=RADER( A10:B12) returnerar 3.  
=RADER( hare) ger 2 om "hare "är det namngivna området (C1:D3).  
Funktionen RADER visar fr o m %PRODUCTNAME 5.0 ett annat tolkningssätt än i tidigare versioner om Du överlämnar en internt genererad matris som parameter.  
När Du laddar äldre %PRODUCTNAME Calc-dokument och har använt sådana parametrar, bör Du tänka på att RADER() i sådana fall nu returnerar andra resultat (inte kolumnernas antal som tidigare, utan radernas).  
KOLUMNER, RAD.  
Kategori Text  
Här förklaras de funktioner som hör till kategorin Text med hjälp av ett exempel.  
De beskrivs nedan.  
ARABISK  
Beräknar värdet på en romersk siffra.  
Värdeområdet måste ligga mellan 0 och 3999.  
Syntax  
ARABISK( text)  
text är texten som visar en romersk siffra.  
Exempel  
Arabisk( "mxiv") ger resultatet 1014  
Arabisk( "mmii") ger resultatet 2002  
ROMERSK.  
BAS  
Omvandlar ett positivt heltal i en text ur talsystemet till den angivna basen.  
Siffrorna 0-9 och bokstäverna A-Z används.  
Syntax  
BAS( tal; roten ur[; minimilängd])  
tal är ett godtyckligt positivt heltal, som ska konverteras.  
roten ur anger talsystemets bas och är ett positivt heltal mellan 2 och 36.  
Detta är en valfri parameter.  
Om parametern överlämnas, fylls en text, som är mindre än den angivna minimilängden, med nollor åt vänster.  
Exempel  
BAS( 17;10;4) ger 0017 i decimalsystemet.  
BAS( 17;10;4) ger 10001 i det binära systemet.  
BAS( 255;16;4) ger 00FF i det hexadecimala talsystemet.  
DECIMAL.  
KOD  
Här visas koden för det första tecknet i en text eller en sträng.  
Syntax  
KOD( text)  
text är den text för vilken det första tecknets kod ska tas fram..  
Exempel  
KOD( "Hieronymus") ger 72, KOD("hieroglyfisk") ger 104.  
Den här koden är inte ASCII-koden, utan den aktuella kodtabellens kod.  
TECKENKOD.  
DECIMAL  
Omvandlar en text med tecken ur ett talsystem till basen rot i ett decimaltal. rot ska ligga i intervallet 2 till 36.  
Inledande blanktecken och tabbtecken ignoreras, och versaler eller gemener i text saknar betydelse.  
Om rot är lika med 16, ignoreras ett inledande x eller X eller 0x eller 0X och ett avslutande h eller H.  
Om rot är lika med 2, ignoreras ett efterföljande b eller B.  
Andra tecken som inte hör till talsystemet genererar ett fel.  
Syntax  
DECIMAL( text; rot)  
text är den text som ska omvandlas.  
För det t.ex. ska gå att skilja ett hexadecimaltal som A1 från referensen till cell A1 är det nödvändigt att du sätter talet inom citationstecken: t.ex. "A1" eller "AFFE ".  
rot anger talsystemets bas och är ett positivt heltal mellan 2 och 36.  
Exempel  
DECIMAL( "17";10) ger 17.  
DECIMAL( "AFFE";16) ger 45054.  
DECIMAL( "0101";2) ger 5.  
BAS.  
VALUTA  
Med denna funktion kan Du omvandla ett godtyckligt decimaltal till ett belopp med valutaangivelse.  
Därutöver avrundas värdet till antalet decimaler.  
I textfältet värde anger Du det rationella tal som ska omvandlas till valutaformat.  
Du kan också ange det antal decimaler som ska anges i valutaformatet i textfältet D.  
Om inget värde anges, visas talet i valutaformat med två decimaler.  
Syntax  
VALUTA( värde; D)  
värde är ett tal, en referens till en cell, som innehåller ett tal eller en formel, som ger ett tal.  
D är antalet siffror efter kommat.  
Exempel  
VALUTA( 255) visar 255,00 €.  
VALUTA( 367,456;2) ger 367,46 €.  
Använd det decimaltecken som är giltigt enligt den aktuella språkvarianten.  
FASTTAL, TEXT, TEXTNUM.  
ERSÄTT  
Om Du vill byta ut en viss del av en sträng mot en annan sträng, anger Du här den text som ska bytas ut, dess position och längd samt textersättningen.  
Med den här funktionen kan Du byta ut både tecken och tal (som automatiskt omvandlas till text).  
Funktionens resultat är alltid en text.  
Om Du vill fortsätta att räkna med ett utbytt tal, måste Du omvandla resultatet till ett tal med funktionen TEXTNUM.  
Om Du anger en text som inte kan tolkas som ett tal och som inte automatiskt kan omvandlas till text ska texten stå inom citattecken.  
Syntax  
ERSÄTT( text, position, längd; textersättning)  
text är den text i vilken en del ska ersättas.  
position är den teckenposition från och med vilken ersättningen ska göras.  
längd är det antal tecken som ska ersättas.  
textersättning är den text som ska sättas in.  
Exempel  
ERSÄTT( 12345,67;1;1;444) returnerar 4442345,67, formaterat som text.  
Det första tecknet ersätts med den kompletta textersättningen.  
RENSA, SÖK, EXTEXT, BYT.UT.  
FASTTAL  
Här kan du bestämma att ett tal ska visas med ett fast antal decimaler och med eller utan tusentalsavgränsare.  
Du kan använda funktionen för att på ett enhetligt sätt formatera en sifferkolumn med ett fast antal decimaler och med eller utan tusentalsavgränsare.  
Syntax  
FASTTAL( tal; Decimaler; Inga tusentalsavgränsare)  
tal är det tal som ska formateras.  
Decimaler är antalet decimaler som ska visas.  
Inga tusentalsavgränsare (valfritt) definierar om tusentalsavgränsare ska sättas.  
Om Inga tusentalsavgränsare är ett tal inte lika med 0 döljs tusentalsavgränsarna.  
Om Inga tusentalsavgränsare är lika med 0 eller utelämnat visas tusentalsavgränsarna från din aktuella språkvariant.  
Exempel  
FASTTAL( 1234567,89;3) returnerar 1.234.567,890.  
FASTTAL( 1234567,89;3;1) returnerar 1234567, 890.  
VALUTA, AVRUNDA, TEXT, TEXTNUM.  
HITTA  
Om Du vill söka igenom en text efter en viss sträng kan Du i fältet söktext ange den sträng som programmet ska söka efter i den text som Du anger i fältet text.  
Du kan även ange sökningens början.  
Söktexten kan vara en enskild bokstav, ett tal, en godtycklig teckenföljd eller ett ord.  
Sökningsfunktionen skiljer mellan versaler och gemener.  
Syntax  
HITTA( söktext; text; position)  
söktext är den text som det ska sökas efter.  
text är den text i vilken sökningen ska ske.  
position (valfri) är den position i texten från och med vilken sökningen ska ske.  
Exempel  
HITTA( 76;998877665544) returnerar 6.  
EXAKT, LÄNGD, SÖK, EXTEXT.  
RENSA  
Om du vill ta bort blanksteg som står framför en sträng, eller vänsterjustera cellinnehåll, anger du den sträng som ska rensas som parameter text.  
Syntax  
RENSA( text)  
text är den text där inledande blanksteg raderas eller cellen vänsterjusteras.  
Exempel  
RENSA( "hej") returnerar hej.  
ERSÄTT, STÄDA, EXTEXT, BYT.UT.  
VERSALER  
Den följd av bokstäver som Du skriver in i textfältet text omvandlas i sin helhet till versaler.  
Syntax  
VERSALER( text)  
text är texten där små bokstäver ska ersättas med stora.  
Exempel  
VERSALER( "God morgon") returnerar GOD MORGON.  
INITIAL, GEMENER.  
INITIAL  
I den bokstavsföljd som Du skriver in i textfältet text omvandlas den första bokstaven efter varje blanktecken till en versal.  
Syntax  
INITIAL( text)  
text är den text i vilken början på varje ord ska ersättas med versaler.  
Exempel  
INITIAL( "sun microsystems") returnerar Sun Microsystems.  
VERSALER, GEMENER.  
EXAKT  
Om Du vill jämföra två strängar med varandra skriver Du in de strängar som ska jämföras i de båda textfälten.  
Om strängarna överensstämmer blir resultatet SANT.  
Kontrollen tar hänsyn till gemener och versaler.  
Syntax  
EXAKT( text_1; text_2)  
text_1 är den första texten för textjämförelsen.  
text_2 är den andra texten för textjämförelsen.  
Exempel  
EXAKT( "Sun microsystems" ;"Sun Microsystems") returnerar FALSKT.  
LÄNGD, SÖK.  
GEMENER  
Den följd av bokstäver som Du skriver in i textfältet text omvandlas i sin helhet till gemener.  
Syntax  
GEMENER( text)  
text är den text i vilken versaler ska ersättas med gemener.  
Exempel  
GEMENER( "Sun") returnerar sun.  
VERSALER, INITIAL.  
VÄNSTER  
Den här funktionen returnerar det första tecknet eller det första antalet tecken i sträng.  
Syntax  
VÄNSTER( text; antal)  
text är den text vars vänstra förled ska bestämmas.  
antal (valfri) är antalet tecken för det vänstra förledet.  
Om parametern saknas returnereras ett tecken.  
Exempel  
VÄNSTER( "stäng av";3) returnerar stä.  
HÖGER, EXTEXT.  
LÄNGD  
Den här funktionen returnerar längden på en sträng.  
Mellanslag räknas med.  
Syntax  
LÄNGD( text)  
text är den text vars längd ska fastställas.  
Exempel  
LÄNGD( "God dag") ger resultatet 7.  
LÄNGD( 12345,67) ger resultatet 8.  
EXAKT, SÖK.  
HÖGER  
Den här funktionen returnerar det sista tecknet eller det sista antalet tecken i en sträng.  
Syntax  
HÖGER( text; antal)  
text är texten vars högra deltext ska bestämmas.  
antal (valfri) är antalet tecken för den högra deltexten.  
Exempel  
HÖGER( "Din buspojke";5) ger resultatet pojke.  
VÄNSTER, EXTEXT.  
ROMERSK  
Omvandlar ett tal till romerska siffror.  
Värdeområdet måste ligga mellan 0 och 3999, lägets värde är begränsat till 0 och 4.  
Syntax  
ROMERSK( tal; läge)  
tal är talet som ska omvandlas till romerska siffror.  
läge (valfritt) anger graden av förenkling.  
Ju högre värde desto mer förenklas de romerska siffrorna.  
Exempel  
ROMERSK( 999) ger resultatet CMXCIX  
ROMERSK( 999;0) ger resultatet CMXCIX  
ROMERSK( 999;1) ger resultatet LMVLIV  
ROMERSK( 999;2) ger resultatet XMIX  
ROMERSK( 999;3) ger resultatet VMIV  
ROMERSK( 999;4) ger resultatet IM  
ARABISK  
SÖK  
Den här funktionen returnerar positionen för en deltext inom en sträng.  
Alternativt kan du definiera sökningens början.  
Söktexten kan vara ett tal eller en valfri teckenföljd.  
Sökningen är inte versalkänslig.  
Syntax  
SÖK( söktext; text; position)  
söktext är den text som det ska sökas efter.  
text är den text i vilken sökningen ska ske.  
position (valfri) är den position i texten från och med vilken sökningen ska ske.  
Exempel  
SÖK( 54;998877665544) ger resultatet 10.  
SÖK( 11;998877665544) ger resultatet #VÄRDE!.  
ERSÄTT, HITTA, EXTEXT, BYT.UT.  
STÄDA  
Alla tecken som inte kan skrivas ut tas bort från strängen.  
Syntax  
STÄDA( text)  
text är den text ur vilken de tecken som inte kan skrivas ut ska tas bort.  
Exempel  
Om du skriver in (ej utskrivbart tecken) Hallå inom citattecken blir resultatet Hallå.  
RENSA, TECKEN.  
T  
Den här funktionen omvandlar ett tal till en tom textsträng.  
Syntax  
T( värde)  
värde är det värde som ska omvandlas.  
Om den refererade cellen innehåller ett tal eller en formel med numeriskt resultat returneras en tom sträng.  
Exempel  
T( 12345) blir till en tom sträng "" om 12345 är formaterat som tal.  
T( "12345") returnerar 12345.  
N, TEXTNUM.  
EXTEXT  
Den här funktionen returnerar en del av texten från en sträng.  
Den bestämmer startpositionen och antalet tecken.  
Syntax  
EXTEXT( text; start; antal)  
text är den text vars delord ska fastställas.  
start är den position från och med vilken delordet ska fastställas.  
antal är antalet tecken för delordet.  
Exempel  
EXTEXT( "Funktionsautopilot";10;4) ger resultatet auto.  
KOD, HITTA, VÄNSTER, HÖGER, SÖK.  
TEXT  
Den här funktionen omvandlar ett tal till en text.  
Textens utseende anger du i den andra parametern.  
Syntax  
TEXT( tal; format)  
tal är det siffervärde som ska omvandlas.  
format är den text som bestämmer formatet. (Avgörande för resultatet här är vilket språk som har angetts i cellformatet.)  
Exempel  
TEXT( 54321 ;"00,00") ger resultatet 54321,00.  
VALUTA, FASTTAL, T, TEXTNUM.  
SAMMANFOGA  
Om Du vill sammanfoga flera texter till en, skriver Du in de enskilda textpassagerna i textfälten.  
Syntax  
SAMMANFOGA( text 1;...;text 30)  
text 1 till text 30 är upp till 30 texter, som kan kopplas samman till en textkedja.  
Exempel  
SAMMANFOGA( "Hej! ""Hur" "mår ""du?") ger resultatet Hej! Hur mår du?  
BYT.UT  
Om du vill byta ut enskilda textdelar mot andra, kan du ange den text, som innehåller textdelen som ska bytas ut, i fältet text.  
I fältet söktext skriver du in den text som ska ersättas av den text som står i fältet textersättning.  
I fältet förekomst kan du ange vid vilken förekomst söktexten ska ersättas.  
Syntax  
BYT.UT( text; söktext; textersättning; förekomst)  
text är den text i vilken deltexter ska bytas ut.  
söktext är den deltext som ska ersättas (flera gånger).  
textersättning är den text som ska ersätta deltexten.  
förekomst (valfri) anger vid vilken förekomst i ordningen av söktexten ersättningen ska göras.  
Om den här parametern saknas ersätts söktexten överallt.  
Exempel  
BYT.UT( "123123123"; "3"; "abc") ger resultatet 12abc12abc12abc.  
BYT.UT( "123123123"; "3"; "abc"; 2) ger resultatet 12312abc123.  
ERSÄTT, RENSA.  
TEXTNUM  
Den här funktionen omvandlar en text till ett tal.  
Syntax  
TEXTNUM( text)  
text är den text som ska omvandlas till ett tal.  
Exempel  
TEXTNUM( "4321") ger resultatet 4321.  
VALUTA, FASTTAL, TEXT.  
REP  
Den här funktionen mångfaldigar en sträng till ett antal kopior.  
Syntax  
REP( text, antal)  
text är texten som ska upprepas.  
antal är antalet upprepningar.  
Resultatet får vara högst 255 tecken långt.  
Exempel  
REP( "God morgon"; 2) ger resultatet God morgonGod morgon.  
TECKEN  
Den här funktionen omvandlar ett tal till ett tecken motsvarande den aktuella kodtabellen.  
Talet kan vara ett två - eller tresiffrigt naturligt tal.  
Syntax  
TECKEN( tal)  
tal är kodvärdet för tecknet.  
Exempel  
TECKEN( 100) ger resultatet d.  
KOD.  
Kategorin Add-in  
Här kan du använda ytterligare add-in-funktioner.  
Add-in-koncept  
En beskrivning av %PRODUCTNAME Calcs add-in-gränssnitt finns också i hjälpen.  
Där finns också en beskrivning av viktiga funktioner och parametrar för ett Shared Library en %PRODUCTNAME Calc-add-in-DLL.  
Medföljande add-ins  
I %PRODUCTNAME ingår exempel för add-in-gränssnittet i %PRODUCTNAME Calc.  
Om du har installerat add-ins finns Shared Libraries DLL:s i {installpath} / program / addin.  
De genererar funktioner, som du hittar i Funktionsautopiloten under kategorin Add-in.  
Analysfunktioner del 1  
Analysfunktioner del 2  
I add-in-mappen finns det dessutom en underordnad mapp med namnet "source".  
Den innehåller källkoden till Shared Libraries DLL-filerna och ger dig som är intresserad av programmering en inblick i funktionssättet för ett addIn-Shared Library en add-in-DLL.  
"Rot*.  
SO DLL "genererar en krypteringsfunktion med namnet ROT13, som bygger på en enkel algoritm.  
Filen "Dfa*.  
SO DLL "tillhandahåller extra datumfunktioner:  
ÄRSKOTTÅR, ANTALÅR, ANTALMÅNADER, DAGARPÅÅRET, DAGARIMÅNADEN, ANTALVECKOR, VECKORPERÅR.  
Funktionerna som du erhåller med "Dfa*.  
SO DLL "kan du bara använda om standardinställningen i %PRODUCTNAME är aktiverad, med 1899-12-30 som nollpunkt för tidsaxeln under Verktyg - Alternativ - Tabelldokument - Beräkna i området Datum.  
Observera att det finns saker som du måste tänka på när du anger datum.  
ÄRSKOTTÅR  
Beräknar om året, då ett datum infaller, är ett skottår.  
Om så är fallet returnerar den här funktionen värdet 1 (SANT), i annat fall 0 (FALSKT).  
Syntax  
ÄRSKOTTÅR( datum)  
datum:  
Beräkningen ska fastställa om det inträffar under ett skottår.  
Exempel  
ÄRSKOTTÅR( 68.02.29) ger resultatet 1.  
ANTALÅR  
Bestämmer antalet år mellan två datum.  
Syntax  
ANTALÅR( Startdatum, Slutdatum, Typ)  
Startdatum:  
Tidigare datum  
Slutdatum:  
Senare datum  
Typ:  
Bestämmer hur skillnaden ska anges.  
Möjliga värden är 0 (intervall) och 1 (i kalenderår).  
ANTALMÅNADER  
Bestämmer antalet månader mellan två datum.  
Syntax  
ANTALMÅNADER( datum_1, datum_2, typ)  
datum_1:  
Tidigare datum  
datum_2:  
Senare datum  
typ:  
Bestämmer hur skillnaden ska anges.  
Möjliga värden är 0 (intervall) och 1 (i kalendermånader).  
ROT13  
Krypterar en teckensträng genom att förskjuta tecknen 13 positioner i alfabetet.  
Efter bokstaven Z börjar funktionen om från alfabetets början igen (rotation).  
Du dekrypterar texten genom att låta krypteringsfunktionen gå igenom koden igen.  
Syntax  
ROT13( text)  
text:  
Anger den teckensträng som ska krypteras.  
ROT13( ROT13(text)) dekrypterar koden igen.  
Exempel  
ROT13( "Detta är en hemlig kod") ger resultatet "Qrggn äe ra urzyvt xbg ".  
ROT13( "Qrggn ine ra urzyvt xbq") ger resultatet "Detta var en hemlig kod ".  
DAGARPÅÅRET  
Bestämmer antalet dagar per år för ett datum.  
Syntax  
DAGARPÅÅRET( datum)  
datum:  
Datum, för vilket antalet dagar per år ska bestämmas.  
Exempel  
DAGARPÅÅRET( 68-02-29) returnerar 366 dagar.  
DAGARIMÅNADEN  
Bestämmer antalet dagar per månad för ett datum.  
Syntax  
DAGARIMÅNADEN( datum)  
datum:  
Datum, för vilket antalet dagar per månad ska bestämmas.  
Exempel  
DAGARIMÅNADEN( 68-02-17) returnerar 29 dagar.  
ANTALVECKOR  
Bestämmer antal veckor mellan två datum.  
Syntax  
ANTALVECKOR( datum_1, datum_2, typ)  
datum_1:  
Tidigare datum  
datum_2:  
Senare datum  
typ:  
Bestämmer hur skillnaden ska anges.  
Möjliga värden är 0 (intervall) och 1 (i kalenderveckor).  
VECKORPERÅR  
Bestämmer antalet veckor per år för ett datum.  
Kalenderveckan definieras så att en kalendervecka vid ett årsskifte räknas till det år där flest dagar i den veckan infaller.  
Syntax  
VECKORPERÅR( datum)  
datum:  
Datum, för vilket antalet veckor per år ska bestämmas.  
Exempel  
VECKORPERÅR( 70-02-17) returnerar 53.  
Add-ins via %PRODUCTNAME API  
Add-ins kan, förutom som DLL, även implementeras via %PRODUCTNAME API.  
Du måste definiera en tjänst som stöder com::sun::star::sheet::AddIn och en implementering av denna måste registreras.  
Ytterligare information, som förutsätter ingående kunskaper om %PRODUCTNAME API-dokumentation, kan erhållas på begäran.  
Programmera Add-in till %PRODUCTNAME Calc  
I %PRODUCTNAME Calc kan du integrera en add-in, d.v.s. en extern programmodul, som ger dig ytterligare funktioner när du arbetar med kalkylprogrammet.  
Dessa visas i Funktionsautopiloten under kategorin Add-in.  
Om du själv vill programmera en sådan add-in-modul, får du här reda på vilka funktioner Shared Library externa DLL:er ska exportera så att add-in-programmet kan integreras ordentligt.  
%PRODUCTNAME letar efter en underordnad mapp, "addin", i den sökväg för moduler som du har angett under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar och söker i denna efter en lämplig Shared Library DLL.  
För att denna DLL ska kunna identifieras av %PRODUCTNAME, måste den ha vissa egenskaper som beskrivs nedan.  
Med hjälp av den här informationen kan du programmera en egen add-in till Funktionsautopiloten i %PRODUCTNAME Calc.  
I programpaketet finns två exempel för add-in-gränssnittet i %PRODUCTNAME Calc.  
Om du angav att även add-ins skulle installeras när du installerade programmet, innehåller Office-mappen en "addin"-mapp som, vid sidan av exempel-DLL:erna, innehåller en ytterligare underordnad mapp, "source", i vilken källkoden finns.  
En beskrivning av de add-in-funktioner som du får genom exempel-DLL:erna hittar du under kategorin Add-in i %PRODUCTNAME Calc-hjälpen till funktionsautopiloten.  
Add-in-konceptet  
Varje add-in-bibliotek innehåller flera funktioner.  
Några av dem är förvaltningsfunktioner som måste uppfylla en viss konvention.  
Med dessa funktioner kan du få information om de övriga funktionerna som utgör den egentliga utökningen av %PRODUCTNAME Calc.  
Namnen på de här funktionerna är godtyckliga, men de måste följa vissa regler vad gäller överlämnandet av parametrar.  
Den exakta namngivningen och anropskonventionerna är plattformsberoende.  
Pascalkonventionerna, eftersom Pascal fortfarande används mycket i Windows-miljön.  
Shared Library Add-in-DLL -funktioner  
I det enklaste fallet ska förvaltningsfunktionerna GetFunctionCount och GetFunctionData finnas.  
Med dessa kan Du bestämma antalet funktioner, parametertyper och returvärden.  
För resultatvärden stöds typerna Double och String.  
Vad gäller parametrar stöds dessutom cellområdena Double Array, String Array och Cell Array.  
Parametrar överlämnas per referens.  
Därför kan du i allmänhet ändra värdena.  
Detta stöds dock inte av %PRODUCTNAME Calc, eftersom det inte är meningsfullt i ett kalkylprogram.  
Du kan ladda bibliotek under körtid och analysera deras innehåll med de båda administrationsfunktionerna.  
För varje funktion ges information om parametrarnas antal och typ, ett programinternt namn, det verkliga namnet och ett administrationsnummer.  
Funktionerna anropas synkront och returnerar omedelbart sina resultat.  
Realtimefunktioner (asynkrona funktioner) är visserligen också möjliga, men de är för komplexa för att närmare förklaras här.  
Allmänt om gränssnittet  
Det maximala antalet parametrar i en AddIn-funktion som integrerats i %PRODUCTNAME Calc är 16: ett resultatvärde och maximalt 15 input-funktionsparametrar.  
Datatyperna är definierade på följande sätt:  
Datatyp  
Definition  
CALLTYPE  
under Windows:  
FAR PASCAL (_far _pascal)  
annars: default (operativsystemsspecifik standard)  
USHORT  
2 byte unsigned Integer  
double  
8 byte plattformsberoende format  
Paramtype  
plattformsberoende som int  
PTR_DOUBLE =0 pekare på en double  
PTR_STRING =1 pekare på en noll-terminerad teckenkedja  
PTR_DOUBLE_ARR =2 pekare på en Double Array  
PTR_DOUBLE_ARR =3 pekare på en String Array  
PTR_DOUBLE_ARR =4 pekare på en Cell Array  
NONE =5  
Shared Library DLL -funktioner  
Nedan beskrivs de funktioner som anropas vid ett Shared Library en extern DLL.  
För alla Shared Library DLL -funktioner gäller:  
void CALLTYPE fn( out, in1, in2,...)  
Output:  
Resultatvärde  
Input:  
Godtyckligt antal valfria typer (double&, char*, double*, char**, Zellbereich), varvid cellområdet är en Array av typen Double Array, String Array eller Cell Array.  
GetFunctionCount()  
Returnerar antalet funktioner utan förvaltningsfunktionerna i referensparametern.  
Varje funktion har ett entydigt nummet mellan 0 och nCount-1.  
Detta nummer används senare för funktionerna GetFunctionData och GetParameterDescription.  
Syntax  
void CALLTYPE GetFunctionCount( USHORT& nCount)  
Parameter  
USHORT &nCount:  
Output:  
Referens till variabel, som ska innehålla antalet AddIn-funktioner.  
Om AddIn-programmet t ex ställer 5 funktioner till %PRODUCTNAME Calcs förfogande är nCount=5.  
GetFunctionData()  
Bestämmer alla viktig information till en AddIn-funktion  
Syntax  
void CALLTYPE GetFunctionData( USHORT& nNo, char* pFuncName, USHORT& nParamCount, Paramtype* peType, char* pInternalName)  
Parameter  
USHORT& nNo:  
Input:  
Funktionsnummer mellan 0 och nCount-1 inklusive.  
char* pFuncName:  
Output:  
Funktionsnamn ur programmerarens synvinkel, så som det betecknas i Shared Library DLL.  
Detta namn bestämmer inte beteckningen i funktionsautopiloten.  
USHORT& nParamCount:  
Output:  
Antal parametrar för AddIn-funktionen.  
Maximivärdet är 16.  
Paramtype* peType:  
Output:  
Pekare på en Array med exakt 16 variabler av typen Paramtype.  
De första nParaCount-posterna fylls med typen för respektive parameter.  
char* pInternalName:  
Output:  
Funktionsnamn ur användarens synvinkel, så som det visas i funktionsautopiloten.  
Kan innehålla omljud.  
Parametrarna pFuncName och pInternalName är char Arrays som implementerats med storleken 256 i %PRODUCTNAME Calc.  
GetParameterDescription()  
Ger en kort beskrivning av AddIn-funktionen och dess parametrar.  
Denna funktion kan Du, om Du vill, använda för att visa en funktions - och parameterbeskrivning.  
Syntax  
void CALLTYPE GetParameterDescription( USHORT& nNo, USHORT& nParam, char* pName, char* pDesc)  
Parameter  
USHORT& nNo:  
Input:  
Funktionens nummer i biblioteket mellan 0 och nCount-1.  
USHORT& nParam:  
Input:  
Parametrar börjar vid 1.  
Om nParam är 0 ska beskrivningen av funktionen i sig ges i pDesc. pName är i detta fall betydelselös.  
char* pName:  
Output:  
Upptar namnet respektive parametertypen, t ex ordet "Tal" eller "Teckenkedja "eller "Datum" eller liknande.  
Implementeras som char[ 256] i %PRODUCTNAME Calc.  
char* pDesc:  
Output:  
Antar parameterns beskrivning, t ex "Värde med vilket universum ska beräknas".  
Implementeras som char[ 256] i %PRODUCTNAME Calc.  
pName och pDesc är char Arrays, som implementerats med storleken 256 i %PRODUCTNAME Calc.  
Tänk på att den plats som står till förfogande i funktionsautopiloten är begränsad och att de 256 tecknen inte kan utnyttjas i sin helhet.  
Cellområden  
I följande tabell ser Du vilka datastrukturer en extern programmodul måste tillhandahålla för att överlämna cellområden. %PRODUCTNAME Calc skiljer mellan tre olika Arrays, beroende på datatyp.  
Double Array  
Du kan överlämna ett cellområde med värden av typen tal / double som parameter.  
En Double Array definieras på följande sätt i %PRODUCTNAME Calc:  
Offset  
Namn  
Beskrivning  
0  
Col1  
Kolumnnummer i cellområdets övre vänstra hörn.  
Räkningen börjar med 0.  
2  
Row1  
Radnummer i cellområdets övre vänstra hörn, räknat från 0.  
4  
Tab1  
Tabellnummer i cellområdets övre vänstra hörn, räknat från 0.  
6  
Col2  
Kolumnnummer i cellområdets nedre högra hörn.  
Räkningen börjar med 0.  
8  
Row2  
Radnummer i cellområdets nedre högra hörn, räknat från 0.  
10  
Tab2  
Tabellnummer i cellområdets nedre högra hörn, räknat från 0.  
12  
Count  
Antal följande element.  
Tomma celler räknas inte och överlämnas inte.  
14  
Col  
Elementets kolumnnummer.  
Räkningen börjar med 0.  
16  
Row  
Elementets radnummer, räknat från 0.  
18  
Tab  
Elementets tabellnummer, räknat från 0.  
20  
Error  
Felnummer, varvid värdet 0 för "inget fel" är belagt.  
När elementet kommer från en formelcell, bestäms felvärdet av formeln.  
22  
Value  
8 byte IEEE-variabel av typen double / flytande komma  
30  
...  
Nästa element  
String Array  
Ett cellområde, som innehåller värden av datatypen Text överlämnas som String Array.  
En String Array definieras på följande sätt i %PRODUCTNAME Calc:  
Offset  
Namn  
Beskrivning  
0  
Col1  
Det övre vänstra hörnets kolumnnummer i cellområdet.  
Räkningen börjar med 0.  
2  
Row1  
Radnummer i cellområdets övre vänstra hörn, räknat från 0.  
4  
Tab1  
Tabellnummer i cellområdets övre vänstra hörn, räknat från 0.  
6  
Col2  
Kolumnnummer i cellområdets nedre högra hörn.  
Räkningen börjar med 0.  
8  
Row2  
Radnummer i cellområdets nedre högra hörn, räknat från 0.  
10  
Tab2  
Tabellnummer i cellområdets nedre högra hörn, räknat från 0.  
12  
Count  
Antal följande element.  
Tomma celler räknas inte och överlämnas inte.  
14  
Col  
Elementets kolumnnummer.  
Räkningen börjar med 0.  
16  
Row  
Elementets radnummer, räknat från 0.  
18  
Tab  
Elementets tabellnummer, räknat från 0.  
20  
Error  
Felnummer, varvid värdet 0 för "inget fel" är belagt.  
När elementet kommer från en formelcell, bestäms felvärdet av formeln.  
22  
Len  
Längden hos den följande strängen, inklusive avslutande noll-byte.  
När längden inklusive avslutande noll-byte ger ett udda värde läggs ytterligare en noll-byte till värdet, så att ett jämnt värde fås.  
Därför beräknas Len med ((StrLen+2)&~1).  
24  
String  
Teckenföljd med avslutande noll-byte.  
24+Len  
...  
Nästa element  
Cell Array  
Använd Cell Arrays om Du vill anropa cellområden som kan innehålla både text och siffror.  
En Cell Array definieras på följande sätt i %PRODUCTNAME Calc:  
Offset  
Namn  
Beskrivning  
0  
Col1  
Det övre vänstra hörnets kolumnnummer i cellområdet.  
Räkningen börjar med 0.  
2  
Row1  
Radnummer i cellområdets övre vänstra hörn, räknat från 0.  
4  
Tab1  
Tabellnummer i cellområdets övre vänstra hörn, räknat från 0.  
6  
Col2  
Kolumnnummer i cellområdets nedre högra hörn.  
Räkningen börjar med 0.  
8  
Row2  
Radnummer i cellområdets nedre högra hörn, räknat från 0.  
10  
Tab2  
Tabellnummer i cellområdets nedre högra hörn, räknat från 0.  
12  
Count  
Antal följande element.  
Tomma celler räknas inte och överlämnas inte.  
14  
Col  
Elementets kolumnnummer.  
Räkningen börjar med 0.  
16  
Row  
Elementets radnummer, räknat från 0.  
18  
Tab  
Elementets tabellnummer, räknat från 0.  
20  
Error  
Felnummer, varvid värdet 0 för "inget fel" är belagt.  
När elementet kommer från en formelcell, bestäms felvärdet av formeln.  
22  
Type  
Cellinnehållets typ, 0 == Double, 1 == String  
24  
Value or Len  
När typ == 0:  
8 byte IEEE-variabel av typen double / flytande komma  
När typ == 1:  
Längden hos den följande strängen, inklusive avslutande noll-byte.  
När längden inklusive avslutande noll-byte ger ett udda värde läggs ytterligare en noll-byte till värdet, så att ett jämnt värde fås.  
Därför beräknas Len med ((StrLen+2)&~1).  
26 if Type==1  
String  
När typ == 1:  
Teckenföljd med avslutande noll-byte.  
32 or 26+Len  
...  
Nästa element  
Kategori Add-in, lista över analysfunktioner del 1  
BESSELI, BESSELJ, BESSELK, BESSELY, BIN.TILL.DEC, BIN.TILL.HEX, BIN.TILL.OKT, DELTA, DEC.TILL.BIN, DEC.TILL.HEX, DEC.TILL.OKT, FELF, FELK, HEX.TILL.BIN, HEX.TILL.DEC, HEX.TILL.OKT, SLSTEG  
Allmän omräkningsfunktion BAS  
Analysfunktioner del 4  
Tillbaka till översiktssidan  
BESSELI  
Här beräknas den modifierade Bessel-funktionen.  
Syntax  
BESSELI( x;n)  
x: värdet som funktionen beräknas för.  
n: ordningstalet för Bessel-funktionen.  
BESSELJ  
Här beräknas Besselfunktionen (cylinderfunktion).  
Syntax  
BESSELJ( x;n)  
x: värdet som funktionen ska beräknas för.  
n: ordningstalet för Bessel-funktionen.  
BESSELK  
Här beräknas den modifierade Bessel-funktionen.  
Syntax  
BESSELK( x;n)  
x: värdet som funktionen beräknas för.  
n: ordningstalet för Bessel-funktionen.  
BESSELY  
Här beräknas den modifierade Bessel-funktionen.  
Syntax  
BESSELY( x;n)  
x: värdet som funktionen beräknas för.  
n: ordningstalet för Bessel-funktionen.  
BIN.TILL.DEC  
Resultatet är det decimala talet av det angivna binära talet.  
Syntax  
BIN.TILL.DEC( Tal)  
Tal: det binära talet.  
Talet får bestå av högst 10 tecken (bitar).  
Den mest signifikanta biten är teckenbiten.  
Negativa tal anges som tvåkomplement.  
Exempel  
=BIN.TILL.DEC( 1100100) ger resultatet 100.  
BIN.TILL.HEX  
Resultatet är det hexadecimala talet av det angivna binära talet.  
Syntax  
BIN.TILL.HEX( Tal;Antal siffror)  
Tal: det binära talet.  
Talet får bestå av högst 10 tecken (bitar).  
Den mest signifikanta biten är teckenbiten.  
Negativa tal anges som tvåkomplement.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=BIN.TILL.HEX( 1100100;6) ger resultatet 000064.  
BIN.TILL.OKT  
Resultatet är det oktala talet av det angivna binära talet.  
Syntax  
BIN.TILL.OKT( Tal;Antal siffror)  
Tal: det binära talet.  
Talet får högst bestå av 10 tecken (bits).  
Den mest signifikanta biten är teckenbiten.  
Negativa tal anges som tvåkomplement.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=BIN.TILL.OKT( 1100100;4) ger resultatet 0144.  
DELTA  
Resultatet är SANT (1) om båda talen som anges som argument är lika annars FALSKT (0).  
Syntax  
DELTA( Tal 1;Tal 2)  
Exempel  
=DELTA( 1;2) ger resultatet 0.  
DEC.TILL.BIN  
Resultatet är det binära talet av det angivna decimala talet mellan -512 och 511.  
Syntax  
DEC.TILL.BIN( Tal;Antal siffror)  
Tal: det decimala talet.  
Om Tal är negativt, returnerar funktionen ett binärt tal som består av 10 tecken.  
Den mest signifikanta biten är teckenbiten, de andra 9 bitarna ger värdet.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=DEC.TILL.BIN( 100;8) ger resultatet 01100100.  
DEC.TILL.HEX  
Resultatet är det hexadecimala talet av det angivna decimala talet.  
Syntax  
DEC.TILL.HEX( Tal;Antal siffror)  
Tal: det decimala talet.  
Om Tal är negativt, returnerar funktionen ett hexadecimalt tal som består av 10 tecken (40 bitar).  
Den mest signifikanta biten är teckenbiten, de andra 39 bitarna ger värdet.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=DEC.TILL.HEX( 100;4) ger resultatet 0064.  
DEC.TILL.OKT  
Resultatet är det oktala talet av det angivna decimala talet.  
Syntax  
DEC.TILL.OKT( Tal;Antal siffror)  
Tal: det decimala talet.  
Om Tal är negativt, returnerar funktionen ett oktalt tal som består av 10 tecken (30 bitar).  
Den mest signifikanta biten är teckenbiten, de andra 29 bitarna ger värdet.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=DEC.TILL.OKT( 100;4) ger resultatet 0144.  
FELF  
Funktionen returnerar värdena från Gauss 'felfunktion.  
Syntax  
FELF( Undre gräns;Övre gräns)  
Undre gräns: integralens undre gräns.  
Övre gräns: valfritt, integralens övre gräns.  
Om det här värdet saknas beräknas mellan 0 och Undre gräns.  
Exempel  
=FELF( 0;1) ger resultatet 0,842701.  
FELFK  
Funktionen returnerar komplementära värden för Gauss 'felfunktion mellan x och oändligt.  
Syntax  
FELFK( Undre gräns)  
Undre gräns: integralens undre gräns.  
Exempel  
=FELFK( 1) ger resultatet 0,157299.  
SLSTEG  
Resultatet är 1 om Tal är större än eller lika med Tröskelvärde.  
Syntax  
SLSTEG( Tal;Tröskelvärde)  
Exempel  
=SLSTEG( 5;1) ger resultatet 1.  
HEX.TILL.BIN  
Resultatet är det binära talet av det angivna hexadecimala talet.  
Syntax  
HEX.TILL.BIN( Tal;Antal siffror)  
Tal: det hexadecimala talet.  
Talet får bestå av högst 10 tecken.  
Den mest signifikanta biten är teckenbiten, de följande bitarna ger värdet.  
Negativa tal anges som tvåkomplement.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=HEX.TILL.BIN( 64;8) ger resultatet 01100100.  
HEX.TILL.DEC  
Resultatet är det decimala talet av det angivna hexadecimala talet.  
Syntax  
HEX.TILL.DEC( Tal)  
Tal: det hexadecimala talet.  
Talet får bestå av högst 10 tecken.  
Den mest signifikanta biten är teckenbiten, de följande bitarna ger värdet.  
Negativa tal anges som tvåkomplement.  
Exempel  
=HEX.TILL.DEC( 64) ger resultatet 100.  
HEX.TILL.OKT  
Resultatet är det oktala talet av det angivna hexadecimala talet.  
Syntax  
HEX.TILL.OKT( Tal;Antal siffror)  
Tal: det hexadecimala talet.  
Talet får bestå av högst 10 tecken.  
Den mest signifikanta biten är teckenbiten, de följande bitarna ger värdet.  
Negativa tal anges som tvåkomplement.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=HEX.TILL.OKT( 64;4) ger resultatet 0144.  
Kategori Add-in, lista över analysfunktioner del 2  
DUBBELFAKULTET, IMARGUMENT, IMABS, IMAGINÄR, IMCOS, IMDIFF, IMDIV, IMEUPPHÖJT, IMKONJUGAT, IMLN, IMLOG10, IMLOG2, IMPRODUKT, IMREAL, IMROT, IMSIN, IMSUM, IMUPPHÖJT, KOMPLEX, KONVERTERA, OKTTILLBIN, OKTTILLDEC, OKTTILLHEX.  
Kategori Statistik  
Analysfunktioner del 1  
Tillbaka till översiktssidan  
IMABS  
Resultatet är absolutvärdet av ett komplext tal.  
Syntax  
IMABS( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMABS( "5+12j") ger resultatet 13.  
IMAGINÄR  
Resultatet är den imaginära andelen av ett komplext tal.  
Syntax  
IMAGINÄR( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMAGINÄR( "4+3j") ger resultatet 3.  
IMUPPHÖJT  
Resultatet är heltalspotensen av ett komplext tal.  
Syntax  
IMUPPHÖJT( Komplext tal;Potens)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Potens: exponenten.  
Exempel  
=IMUPPHÖJT( "2+3i";2) ger resultatet -5+12i.  
IMARGUMENT  
Resultatet är argumentet (vinkeln phi) av ett komplext tal.  
Syntax  
IMARGUMENT( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMARGUMENT( "3+4j") ger resultatet 0,927295.  
IMCOS  
Resultatet är cosinus av ett komplext tal.  
Syntax  
IMCOS( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMCOS( "3+4j") ger resultatet -27.03-3.85i (avrundat).  
IMDIV  
Resultatet är divisionen av två komplexa tal.  
Syntax  
IMDIV( Täljare;Nämnare)  
Täljare, Nämnare: de komplexa talen anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMDIV( "-238+240i" ;"10+24i") ger resultatet 5+12i.  
IMEUPPHÖJT  
Resultatet är e (det Eulerska talet) upphöjt till det komplexa talet.  
Syntax  
IMEUPPHÖJT (Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMEUPPHÖJT ("1+j") ger resultatet 1.47+2.29j (avrundat).  
IMKONJUGAT  
Resultatet är det konjugerade komplexa komplementet till ett komplext tal.  
Syntax  
IMKONJUGAT( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMKONJUGAT( "1+j") ger resultatet 1-j.  
IMLN  
Resultatet är den naturliga logaritmen för ett komplext tal.  
Syntax  
IMLN( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMLN( "1+j") ger resultatet 0.35+0.79j (avrundat).  
IMLOG10  
Resultatet är 10-logaritmen för ett komplext tal.  
Syntax  
IMLOG10( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMLOG10( "1+j") ger resultatet 0.15+0.34j (avrundat).  
IMLOG2  
Resultatet är 2-logaritmen av ett komplext tal.  
Syntax  
IMLOG2( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMLOG2( "1+j") ger resultatet 0.50+1.13j (avrundat).  
IMPRODUKT  
Resultatet är produkten av upp till 29 komplexa tal.  
Syntax  
IMPRODUKT( Komplext tal;Komplext tal 1;...)  
Komplext tal: de komplexa talen anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMPRODUKT( "3+4j" ;"5-3j") ger resultatet 27+11j.  
IMREAL  
Resultatet är realkoefficienten av ett komplext tal.  
Syntax  
IMREAL( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMREAL( "1+3j") ger resultatet 1.  
IMSIN  
Resultatet är sinus av ett komplext tal.  
Syntax  
IMSIN( Komplext tal)  
Komplext tal: det komplexa talet anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMSIN( "3+4j") ger resultatet 3.85+27.02j (avrundat).  
IMDIFF  
Resultatet är subtraktionen av två komplexa tal.  
Syntax  
IMDIFF( Komplext tal 1;Komplext tal 2)  
Komplext tal: de komplexa talen anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMDIFF( "13+4j" ;"5+3j") ger resultatet 8+j.  
IMSUM  
Resultatet är summan av upp till 29 komplexa tal.  
Syntax  
IMSUM( Komplext tal 1;Komplext tal 2;...)  
Komplext tal: de komplexa talen anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMSUM( "13+4j" ;"5+3j") ger resultatet 18+7j.  
IMROT  
Resultatet är roten av ett komplext tal.  
Syntax  
IMROT( Komplext tal)  
Komplext tal: de komplexa talen anges enligt mönstret "x + yi" eller "x + yj ".  
Exempel  
=IMROT( "3+4i") ger resultatet 2+1i.  
KOMPLEX  
Resultatet är ett komplext tal som returneras av realdel och imaginärdel.  
Syntax  
KOMPLEX( Realdel;Imaginärdel;Suffix)  
Realdel: realdelen till det komplexa talet.  
Imaginärdel: imaginärdelen till det komplexa talet.  
Suffix: valfritt, "i" eller "j ".  
Exempel  
=KOMPLEX( 3;4;j) ger resultatet 3+4j.  
OKT.TILL.BIN  
Resultatet är det binära talet av det angivna oktala talet.  
Syntax  
OKT.TILL.BIN( Tal;Antal siffror)  
Tal: det oktala talet.  
Talet får bestå av högst 10 tecken.  
Den mest signifikanta biten är teckenbiten, de följande bitarna ger värdet.  
Negativa tal anges som tvåkomplement.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=OKT.TILL.BIN( 3;3) ger resultatet 011.  
OKT.TILL.DEC  
Resultatet är det decimala talet av det angivna oktala talet.  
Syntax  
OKT.TILL.DEC( Tal)  
Tal: det oktala talet.  
Talet får bestå av högst 10 tecken.  
Den mest signifikanta biten är teckenbiten, de följande bitarna ger värdet.  
Negativa tal anges som tvåkomplement.  
Exempel  
=OKT.TILL.DEC( 144) ger resultatet 100.  
OKT.TILL.HEX  
Resultatet är det hexadecimala talet av det angivna oktala talet.  
Syntax  
OKT.TILL.HEX( Tal;Antal siffror)  
Tal: det oktala talet.  
Talet får bestå av högst 10 tecken.  
Den mest signifikanta biten är teckenbiten, de följande bitarna ger värdet.  
Negativa tal anges som tvåkomplement.  
Antal siffror: antalet siffror som ska användas.  
Exempel  
=OKT.TILL.HEX( 144;4) ger resultatet 0064.  
KONVERTERA_ADD  
Omvandlar ett värde från en måttenhet till motsvarande värde i en annan måttenhet.  
Måttenheterna anger du direkt som text med citattecken eller som referens.  
Om du matar in måttenheterna i celler måste skrivsättet (stor och liten bokstav) överensstämma exakt med följande lista.  
Om du t.ex. vill mata in den lilla bokstaven l (för liter) i en cell matar du in apostrof 'direkt följt av ett l.  
Egenskap  
Enheter  
Massa  
g, sg, lbm, u, ozm, stone, ton, grain, pweight, hweight, shweight  
Längd  
m, mi, Nmi, in, ft, yd, ang, Pica, ell, parsec  
Tid  
yr, day, hr, mn, sec  
Tryck  
Pa, atm, mmHg, torr, psi  
Kraft  
N, dyn, pond  
Energi  
J, e, c, cal, eV, HPh, Wh, BTU  
Effekt  
W, HP, hk  
Magnetism  
T, ga  
Temperatur  
C, F, K, Reau, Rank  
Volym  
l, tsp, tbs, oz, cup, pt, qt, gal, m3, mi3, Nmi3, in3, ft3, yd3, ang3, Pica3, barrel, bushel, regton, Schooner, Middy, Glass  
Yta  
m2, mi2, Nmi2, in2, ft2, yd2, ang2, Pica2, Morgen, ar, acre, ha  
Hastighet  
m / s, m / h, mph, kn, admkn  
Det får stå ett prefixtecken framför varje måttenhet från följande lista:  
Tillåtna prefixtecken  
10^( <0)  
d, c, m, u, n, p, f, a, z, y  
10^( >0)  
e, h, k, M, G, T, P, E, Z, Y  
Syntax  
KONVERTERA_ADD( Tal;Ursprungsenhet;Ny enhet)  
Tal: talet som räknas om.  
Ursprungsenhet: måttenheten för talet som räknas om.  
Ny enhet: måttenheten som talet räknas om till.  
Exempel  
=KONVERTERA_ADD( 10 ;"HP" ;"HK") ger avrundat till två decimaler resultatet 10,14.  
10 hp är 10,14 hk.  
=KONVERTERA_ADD( 10 ;"km" ;"mi") ger avrundat till två decimaler resultatet 6,21.  
K:et är det tillåtna prefixtecknet för faktorn 10^3.  
DUBBELFAKULTET  
Resultatet är fakulteten för talet med steglängd 2.  
Syntax  
DUBBELFAKULTET( Tal)  
Tal: om tal är jämnt beräknas följande fakultet: n*( N-2)*(n-4 )*...*4*2.  
om tal är udda beräknas följande fakultet: n*( N-2)*(n-4 )*...*3*1.  
Exempel  
DUBBELFAKULTET( 6) ger resultatet 48.  
Kategori Finans del 3  
Till finansfunktionerna del 1  
Till finansfunktionerna del 2  
FÖRRÄNTNING, KUPANT, KUPDAGB, KUPDAGBB, KUPDAGNK, KUPFKD, KUPNKD, PERIODER RBETALNING, RRI, RÄNTA, SLUTVÄRDE, UDDAFAVKASTNING, UDDAFPRIS, UDDASAVKASTNING, UDDASPRIS, VDEGRAVSKR, XIRR, XNUVÄRDE, ÅRSRÄNTA.  
UDDAFPRIS  
Beräknar kursen per 100 valutaenheter nominellt värde för ett värdepapper om det första kupongdatumet infaller oregelbundet.  
Syntax  
UDDAFPRIS( Betalning;Förfallodag;Emission; Första kupongdatum;Ränta;Avkastning;Inlösningsvärde;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Emission: datum för värdepappersemissionen.  
Första kupongdatum: värdepapperets första räntedatum.  
Ränta: den årliga räntesatsen.  
Avkastning: den årliga avkastningen på värdepapperet.  
Inlösningsvärde: inlösningsvärdet per 100 valutaenheter nominellt värde.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Betalning:  
11 november 1999, Förfallodag:  
1 mars 2012, Emission:  
15 oktober 1999; Första kupongdatum:  
1 mars 2000.  
Ränta:  
7,85 procent, Avkastning:  
6,25 procent, Inlösningsvärde:  
100 valutaenheter, betalningarnas Frekvens: halvårsvis = 2, Bas: = 1  
Kursen per 100 valutaenheter nominellt värde för ett värdepapper som har ett oregelbundet första räntedatum, beräknas på följande sätt:  
=UDDAFPRIS( "1999-11-11" ;"2012-03-01" ;"1999-10-15" ;"2000-03-01";0,0785;0,0625;100;2;1) returnerar 113,5985  
UDDAFAVKASTNING  
Beräknar avkastningen på ett värdepapper om det första kupongdatumet infaller oregelbundet.  
Syntax  
UDDAFAVKASTNING( Betalning;Förfallodag;Emission; Första kupongdatum;Ränta;Pris;Inlösningsvärde; Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Emission: datum för värdepappersemissionen.  
Första kupongdatum: värdepapperets första räntedatum.  
Ränta: den årliga räntesatsen.  
Pris: värdepapperets pris.  
Inlösningsvärde: inlösningsvärdet per 100 valutaenheter nominellt värde.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Betalning:  
25 januari 1999, Förfallodag:  
1 januari 2004, Emission:  
18 januari 1999; Första kupongdatum:  
15 juli 1999.  
Ränta:  
5,75 procent, Pris:  
84,50 valutaenheter, Inlösningsvärde:  
100 valutaenheter, betalningarnas Frekvens: halvårsvis = 2, Bas: = 0  
Avkastningen på värdepapperet, som har ett oregelbundet första kupongdatum, beräknas på följande sätt:  
=UDDAFAVKASTNING( "1999-01-25" ;"2004-01-01"; "1999-01-18" ;"1999-07-15";0,0575; 84,50; 100;2;0) returnerar 0,097581 eller 9,76%.  
UDDASPRIS  
Beräknar priset per 100 valutaenheter nominellt värde för ett värdepapper om det sista kupongdatumet infaller oregelbundet.  
Syntax  
UDDASPRIS( Betalning;Förfallodag; Sista kupongdatum;Ränta;Avkastning;Inlösningsvärde;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Sista kupongdatum: värdepapperets sista kupongdatum.  
Ränta: den årliga räntesatsen.  
Avkastning: den årliga avkastningen på ett värdepapper.  
Inlösningsvärde: inlösningsvärdet per 100 valutaenheter nominellt värde.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Betalning:  
7 februari 1999, Förfallodag:  
15 juni 1999, Sista kupongdatum:  
15 oktober 1998.  
Ränta:  
3,75 procent, Avkastning:  
4,05 procent, Inlösningsvärde:  
100 valutaenheter, betalningarnas Frekvens: halvårsvis = 2, Bas: = 0  
Priset per 100 valutaenheter nominellt värde för ett värdepapper, som har ett oregelbundet sista kupongdatum, beräknas på följande sätt:  
UDDASPRIS( "1999-02-07" ;"1999-06-15" ;"1998-10-15"; 0,0375; 0,0405;100;2;0) returnerar 99,87829.  
UDDASAVKASTNING  
Beräknar avkastningen på ett värdepapper om det sista kupongdatumet ligger oregelbundet.  
Syntax  
UDDASAVKASTNING( Betalning;Förfallodag; Sista kupongdatum;Ränta;Pris;Inlösningsvärde;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Sista kupongdatum: det sista kupongdatumet för värdepapperet.  
Ränta: den årliga räntesatsen.  
Pris: värdepapperets pris.  
Inlösningsvärde: inlösningsvärdet per 100 valutaenheter nominellt värde.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Betalning:  
20 april 1999, Förfallodag:  
15 juni 1999, Sista kupongdatum:  
15 oktober 1998.  
Ränta:  
3,75 procent, Pris:  
99,875 valutaenheter, Inlösningsvärde:  
100 valutaenheter, betalningarnas Frekvens: halvårsvis = 2, Bas: = 0  
Avkastningen på värdepapperet, som har ett oregelbundet sista kupongdatum, beräknas på följande sätt:  
=UDDASAVKASTNING( "1999-04-20" ;"1999-06-15"; "1998-10-15"; 0,0375; 99,875; 100;2;0) returnerar 0,044873 eller 4,4873%.  
VDB  
Beräknar den artitmetisk-degressiva avskrivningen för en viss period.  
Syntax  
VDEGRAVSKR( AV;RV;LL;Start;Slut;FA;typ)  
AV är tillgångens anskaffningsvärde.  
RV är tillgångens restvärde vid livslängdens slut.  
LL är livslängden uttryckt i antalet avskrivningsperioder.  
S är avskrivningens startperiod.  
Den måste anges i samma tidsenhet som livslängden.  
S är avskrivningens slutperiod.  
FA (valfri) är avskrivningsfaktorn.  
FA=2 betyder dubbel avskrivning.  
Vid typ=0 görs inget byte.  
Exempel  
Hur stor är den aritmetisk-degressiva dubbla avskrivningen för en viss periodiserad tidsrymd, om anskaffningsvärdet är 35 000 valutaenheter och restvärdet 7 500 valutaenheter?  
Livslängden är 3 år.  
Avskrivningen ska beräknas fr.o.m. den 10:e t.o.m. den 20:e perioden.  
VDEGRAVSKR( 35000;7500;36;10;20;2) = 8603,80 valutaenheter.  
Avskrivningen i tidsperioden mellan den 10:e och den 20:e perioden uppgår till 8 603,80 valutaenheter.  
ÅRSAVSKR, DEGAVSKR, LINAVSKR.  
XIRR  
Beräknar internräntan för en lista med betalningar som sker vid olika tidpunkter.  
Om betalningarna görs med jämna mellanrum använder du funktionen IR.  
Syntax  
XIRR( Värden;Tidpunkter;Gissning)  
Värden och tidpunkter: en serie betalningar och de tillhörande datumvärdena.  
Det första dataparet definierar början på betalningsplanen.  
Alla andra datumvärden måste ligga senare men behöver inte vara ordnade.  
Värdeserien måste innehålla minst ett negativt och ett positivt värde (utbetalningar och inbetalningar).  
Gissning: en gissning kan anges för internräntan (valfritt).  
Standard är 10%.  
Exempel  
Beräkna internräntan för följande fem betalningar:  
A  
B  
C  
1  
01-01-01  
-10000  
Utbetalning  
2  
2001-02-01  
2000  
Inbetalningar  
3  
2001-03-15  
2500  
4  
2001-05-12  
5000  
5  
2001-08-10  
1000  
=XIRR( B1:B5; A1:A5; 0,1) returnerar 0,1828.  
XNUVÄRDE  
Beräknar kapitalvärdet (nettonuvärdet) för en lista med betalningar som sker vid olika tidpunkter.  
Om betalningarna sker med jämna mellanrum använder du funktionen NETNUVÄRDE.  
Syntax  
XNUVÄRDE( Ränta;Värden;Tidpunkter)  
Ränta: räntan för betalningarna.  
Värden och tidpunkter: en serie betalningar och tillhörande datumvärden.  
Det första dataparet definierar början på betalningsplanen.  
Alla andra datumvärden måste ligga senare, men behöver inte vara ordnade.  
Värdeserien måste innehålla minst ett negativt och ett positivt värde (utbetalningar och inbetalningar).  
Exempel  
Beräkna kapitalvärdet för de ovannämnda fem betalningarna vid en diskonteringsränta på 6%:  
=XNUVÄRDE( 0,06; B1:B5; A1:A5) returnerar 323,02.  
RRI  
Den här räntefunktionen beräknar räntesatsen som utgör vinsten (avkastningen) på en investering.  
Syntax:  
RRI( P;NUVÄRDE;Slutvärde)  
P är det antal perioder som krävs för beräkningen av räntesatsen.  
Nuvärde är det nuvarande värdet.  
Nuvärdet utgörs av ett insatt belopp eller en naturaförmån av motsvarande värde.  
Du måste ange ett positivt belopp som investering; det får inte vara 0.  
Slutvärde är det värde som investeringen ska uppnå.  
Exempel  
Under en tidsrymd av 4 perioder (år) och med ett nuvärde på 7 000 valutaenheter ska avkastningens räntesats beräknas, när det framtida värdet ska uppgå till 10 000 valutaenheter.  
RRI( 4;7500;10000) = 7,46%  
Förräntningen måste uppgå till 7,46% för att 7 500 valutaenheter ska bli 10 000 valutaenheter.  
LÖPTID.  
RÄNTA  
Beräknar den konstanta räntesatsen för en investering vid regelbundna betalningar.  
Syntax  
RÄNTA( Perioder;Betalning;Nuvärde;Slutvärde;F;gissning)  
Perioder är betalningstiden angiven i antalet perioder.  
Betalning är den konstanta annuiteten som betalas varje period.  
Nuvärde är det nuvarande värdet av varje betalning.  
Slutvärde (valfritt) är det framtida värde som ska ha uppnåtts när alla betalningar är gjorda.  
F = 1 om betalningen görs under periodens början; F = 0 (standardvärde) om den görs vid dess slut.  
gissning (valfritt) är det uppskattade värdet av räntan för den iterativa beräkningen.  
Exempel  
Hur stor är den konstanta räntesatsen vid en betalningstidsrymd på 3 perioder, om 50 valutaenheter betalas regelbundet och nuvärdet är 900 valutaenheter?  
RÄNTA( 3;10;900) = -121%.  
Räntesatsen uppgår alltså till 121%.  
NUVÄRDE, AMORT, BETALNING, RBETALNING, SLUTVÄRDE, PERIODER.  
ÅRSRÄNTA  
Beräknar den årliga räntesatsen som blir resulatet när ett värdepapper (eller annat objekt) köps till ett investeringsvärde och säljs till ett inlösningsvärde.  
Inga räntor betalas.  
Syntax  
ÅRSRÄNTA( Betalning;Förfallodag;Investering;Inlösningsvärde;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet säljs.  
Investering: köppriset.  
Inlösningsvärde: försäljningspriset.  
Exempel  
En tavla köps den 15 januari 1990 för 1 miljon och säljs den 5 maj 2002 för 2 miljoner.  
Hur hög är den genomsnittliga årsräntan?  
=ÅRSRÄNTA( "1990-01-15"; "2002-05-05"; 1000000; 2000000; 3) returnerar 8,12%.  
KUPNKD  
Returnerar den första kupongdagens datum efter likviddagen.  
Formatera resultatet som datum.  
Syntax  
KUPNKD( Betalning;Förfallodag;Frekvens;Bas)  
Betalning: datumet för värdepappersköpet.  
Förfallodag: datumet då värdepapperet förfaller.  
Frekvens: antal räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 25 januari 2001; förfallodagen är den 15 november 2001.  
Räntorna betalas halvårsvis (frekvens är 2).  
När är nästa kupongdatum vid faktisk / 365 beräkning (bas 3)?  
=KUPNKD( "2001-01-25"; "2001-11-15"; 2; 3) ger resultatet 2001-05-15.  
KUPDAGB  
Returnerar antalet dagar i den aktuella ränteperioden i vilken likviddagen ligger som resultat.  
Syntax  
KUPDAGB( Betalning;Förfallodag;Frekvens;Bas)  
Betalning: datumet för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Räntorna betalas halvårsvis (frekvens är 2).  
Hur många dagar finns det i ränteperioden i vilken likviddagen ligger vid faktisk / 365 beräkning (bas 3)?  
=KUPDAGB( "2001-01-25"; "2001-11-15"; 2; 3) ger resultatet 181.  
KUPDAGNK  
Ger antalet dagar från likviddatum till nästa kupongdatum som resultat.  
Syntax  
KUPDAGNK( Betalning;Förfallodag;Frekvens;Bas)  
Betalning: datumet för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 25 januari 2001; förfallodagen är den 15 november 2001.  
Räntorna betalas halvårsvis (frekvens är 2).  
Hur många dagar är det till nästa räntebetalning vid faktisk / 365 beräkning (bas 3)?  
=KUPDAGNK( "2001-01-25"; "2001-11-15"; 2; 3) ger resultatet 110.  
KUPDAGBB  
Returnerar antalet dagar från räntebetalningens första dag för ett värdepapper till likkviddagen.  
Syntax  
KUPDAGBB( Betalning;Förfallodag;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 25 januari 2001; förfallodagen är den 15 november 2001.  
Hur många dagar finns det vid faktisk / 365 beräkning (bas 3)?  
=KUPDAGBB( "2001-01-25"; "2001-11-15"; 2; 3) ger resultatet 71.  
KUPFKD  
Returnerar senaste kupongdatum före likviddagen.  
Formatera resultatet som datum.  
Syntax  
KUPFKD( Betalning;Förfallodag;Frekvens;Bas)  
Betalning: datumet för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Frekvens: antal räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 25 januari 2001; förfallodagen är den 15 november 2001.  
Räntorna betalas halvårsvis (frekvens är 2).  
När var senaste kupongdatum före köpet vid faktisk / 365 beräkning (bas 3)?  
=KUPFKD( "2001-01-25"; "2001-11-15"; 2; 3) returnerar 2000-11-15.  
KUPANT  
Returnerar antalet kuponger (räntebetalningar) mellan likviddatum och förfallodatum.  
Syntax  
KUPANT( Betalning;Förfallodag;Frekvens;Bas)  
Betalning: datumet för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Frekvens: antal räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 25 januari 2001; förfallodagen är den 15 november 2001.  
Hur många kupongdatum finns det vid faktisk / 365 beräkning (bas 3)?  
=KUPANT( "2001-01-25"; "2001-11-15"; 2; 3) returnerar 2.  
RBETALNING  
Beräknar räntan under en period för en investering vid regelbundna betalningar och konstant räntesats.  
Syntax  
RBETALNING( ränta;P;Perioder;Nuvärde;Slutvärde;F)  
ränta är räntesatsen för en periods betalning.  
P är den period för vilken ränta på ränta ska beräknas.  
P=BETALNING om räntan på räntan ska beräknas för den sista perioden.  
Perioder är betalningstiden angiven i antal perioder.  
Nuvärde är det nuvarande värdet av varje betalning.  
Slutvärde (valfritt) är det slutliga värde (framtida värde) som ska ha uppnåtts när alla betalningar är gjorda.  
F = 1 om betalningen görs under periodens början; F = 0 (standardvärde) om den görs vid dess slut.  
Exempel  
Hur stor är förräntningen under den femte perioden (året), om den konstanta räntan är 5% och nuvärdet är 15 000 valutaenheter?  
Den periodiska betalningstiden är sju år.  
RBETALNING( 5%;5;7;15000) = -352,97 valutaenheter.  
Räntan på räntan under den femte perioden (året) uppgår till 352,97 valutaenheter.  
NUVÄRDE, AMORT, KUMRÄNTA, BETALNING, RÄNTA.  
SLUTVÄRDE  
Beräknar slutvärdet av en investering vid regelbundna betalningar och konstant ränta.  
Syntax  
SLUTVÄRDE( ränta; Perioder; Betalning; Nuvärde; F)  
ränta är räntesatsen för en periods betalning.  
Perioder är betalningstiden angiven i antalet perioder.  
Betalning är betalningen för en period.  
Nuvärde (valfritt) är det nuvarande värdet av en investering.  
F (valfritt) definierar förfallotidpunkten för betalningen i början eller i slutet av en period.  
Exempel  
Hur stort är slutvärdet av en investering, om räntesatsen är 4% och betalningstiden vid en periodisk betalning om 750 valutaenheter sträcker sig över två år?  
Investeringens nuvärde är 2 500 valutaenheter.  
Slutvärde( 4%;2;750;2500) = -4234,00 valutaenheter.  
Investeringens slutliga värde är 4 234,00 valutaenheter.  
NUVÄRDE, AMORT, BETALNING, RÄNTA, RBETALNING, PERIODER.  
FÖRRÄNTNING  
Beräknar ett framtida värde av ett begynnelsekapital för en rad periodiskt olika räntesatser.  
Syntax  
FÖRRÄNTNING (Kapital;Räntor)  
Kapital: begynnelsekapital.  
Räntor: en rad räntesatser, t.ex. som område H3:H5 eller som {Lista} (se exempel).  
Exempel  
1000 valutaenheter har placerats på tre år.  
Hur högt är värdet efter tre år?  
=FÖRRÄNTNING( 1000; {0,03; 0,04; 0,05}) returnerar 1124,76.  
PERIODER  
Beräknar antalet betalningsperioder för en investering vid regelbundna betalningar och konstant räntesats.  
Syntax  
PERIODER( ränta;Betalning;Nuvärde;Slutvärde;F)  
ränta är räntesatsen för en periods betalning.  
Betalning är den konstanta annuiteten som ska betalas varje period.  
Nuvärde är det nuvarande värdet av betalningarna.  
Slutvärde (valfritt) är det framtida värde som ska ha uppnåtts när alla betalningar är gjorda.  
F = 1 om betalningen görs under periodens början; F = 0 (standardvärde) om den görs vid dess slut.  
Exempel  
Hur många betalningsperioder omfattar en betalningstid vid en periodisk räntesats på 6%, en periodisk betalning på 153,75 valutaenheter och ett nuvärde på 2 600 valutaenheter?  
PERIODER( 6%;153,75;2600) = -12,02.  
Betalningstidsrymden är alltså 12,02 perioder.  
NUVÄRDE, AMORT, BETALNING, RÄNTA, RBETALNING, SLUTVÄRDE.  
Till finansfunktionerna del 1  
Till finansfunktionerna del 2  
Kategori Finans del 2  
Till finansfunktionerna del 1  
Till finansfunktionerna del 3  
AMORT, BETALNING, BRÅK, DECTAL, KUMPRIS, KUMPRIS_ADD, KUMRÄNTA, KUMRÄNTA_ADD, LINAVSKR, LÖPTID, MLÖPTID, MODIR, NETNUVÄRDE, NOMAVK, NOMAVKDISK, NOMAVKFÖRF, NOMRÄNTA, NOMRÄNTA_ADD, PRIS, PRISDISK, PRISFÖRF, SSVXEKV, SSVXPRIS, SSVXRÄNTA.  
AMORT  
Beräknar den periodiska amorteringen för en investering vid regelbundna betalningar och konstant räntesats.  
Syntax  
AMORT( ränta;P;Perioder;Nuvärde;Slutvärde;F)  
ränta är räntesatsen för en periods betalning.  
P är amorteringsperioden.  
P=1 för den första perioden och P=Perioder för den sista.  
Perioder är betalningstiden angiven i antalet perioder.  
Nuvärde är det nuvarande värdet av varje betalning.  
Slutvärde (valfritt) är det eftersträvade (framtida) värdet.  
F (valfritt) är förfallotidpunkten.  
F = 1 om betalningen görs under periodens början; F = 0 (standardvärde) om den görs vid dess slut.  
Exempel  
Hur hög är den periodiska amorteringen vid en räntesats på 8,75% och en betalningsperiod på 3 år?  
Det nuvarande värdet uppgår till 5.000 valutaenheter.  
Betalning ska alltid göras i början av perioden.  
Det slutliga värdet uppgår till 8.000 valutaenheter.  
AMORT( 8,75%;1;36;5000;8000;1) = -455,98 valutaenheter.  
NUVÄRDE, BETALNING, RÄNTA, RBETALNING, SLUTVÄRDE, PERIODER.  
KUMPRIS  
Beräknar totalbeloppet av amorteringarna för en investering under en viss tidsrymd vid konstant räntesats.  
Syntax  
KUMPRIS( ränta;Perioder;Nuvärde;Start;Slut;F)  
ränta är räntesatsen för en periods betalning.  
Perioder är betalningstiden angiven i antalet perioder.  
Det behöver inte vara ett heltal.  
Nuvärde är det nuvarande värdet av varje betalning.  
Start är den första perioden (startperioden).  
Slut är den sista perioden (slutperioden).  
F = 1 om betalningen görs i periodens början; F = 0 (standardvärde) om den görs i dess slut.  
Exempel  
Hur stor är amorteringsdelen vid 36 perioder och en räntesats på 5,5%?  
Kontantvärdet är 15 000 valutaenheter.  
Amorteringsdelen ska beräknas för en tidsrymd mellan den 10:e och 18:e perioden.  
Förfallodagen är i slutet av perioden.  
KUMPRIS( 5,5%;36;15000;10;18;0) = -2 560,52 valutaenheter.  
Amorteringsandelen mellan den 10:e och 18:e perioden är 2 560,52 valutaenheter.  
KUMRÄNTA.  
KUMPRIS_ADD  
Beräknar den ackumulerade amorteringen på ett lån under en period.  
Syntax  
KUMPRIS_ADD( Ränta;Perioder;Nuvärde;Start;Slut;F)  
Ränta: räntesatsen per period.  
Perioder: totalt antal betalningsperioder.  
Ränta och Perioder måste anges i samma enhet, d.v.s. båda beräknas årsvis eller månadsvis.  
Nuvärde: nuvärdet.  
Startperiod: den första betalningsperioden för beräkningen.  
Slutperiod: den sista betalningsperioden för beräkningen.  
F: förfallotidpunkten för en betalning i slutet av perioden (Typ = 0) eller i början av perioden (Typ = 1).  
Exempel  
Följande hypotekslån tas för ett hus:  
Ränta:  
9,00 procent per år (9% / 12 = 0,0075), löptid:  
30 år (betalningsperioder = 30 * 12 = 360), nuvärde:  
125 000 valutaenheter.  
Hur hög är amorteringen som du betalar det andra året (d.v.s. i perioderna 13 till 24)?  
KUMPRIS_ADD( 0,0075;360;125000;13;24;0) returnerar -934,1071  
Den första månaden betalar du följande amortering:  
KUMPRIS_ADD( 0,0075;360;125000;1;1;0) returnerar -68,27827  
KUMRÄNTA  
Beräknar kumulerade räntor på räntor, d.v.s. totalbeloppet av alla räntor för en investering under en viss tidsperiod.  
Räntesatsen är konstant.  
Syntax  
KUMRÄNTA( ränta;Perioder;Nuvärde;Start;Slut;F)  
Ränta är räntesatsen för en periods betalning.  
Perioder är betalningstiden angiven i antalet perioder.  
Den behöver inte vara ett heltal.  
Nuvärde är det nuvarande värdet av varje betalning.  
Start är den första perioden.  
Slut är den sista perioden.  
F = 1 om betalningen görs i periodens början; F = 0 (standardvärde) om den görs i dess slut.  
Exempel  
Hur stor blir ränteandelen vid en periodisk räntesats på 5,5%, en periodisk tidrymd på 2 år och ett nuvärde på 5 000 valutaenheter?  
Beräkningsperioden börjar med den 4:e och slutar med den 6:e perioden.  
Den periodiska betalningen förfaller i början av perioden.  
KUMRÄNTA( 5,5%;24;5000;4;6;1) = -710,21 valutaenheter.  
Ränteandelen under den 4:e till den 6:e perioden uppgår till 710,21 valutaenheter.  
KUMPRIS  
KUMRÄNTA_ADD  
Beräknar den ackumulerade räntan i en period.  
Syntax  
KUMRÄNTA_ADD( Ränta;Perioder;NUVÄRDE;Startperiod;Slutperiod;Typ)  
Ränta: räntesatsen per period.  
Perioder: totalt antal betalningsperioder.  
Ränta och Perioder måste anges i samma enhet, d.v.s. beräknas årsvis eller månadsvis.  
Nuvärde: nuvärdet.  
Startperiod: den första betalningsperioden för beräkningen.  
Slutperiod: den sista betalningsperioden för beräkningen.  
Typ: förfallotidpunkt för en betalning i slutet av perioden (Typ = 0) eller i början av perioden (Typ = 1).  
Exempel  
Följande hypotekslån tas för ett hus:  
Ränta:  
9,00 procent per år (9% / 12 = 0,0075), löptid:  
30 år (perioder = 30 * 12 = 360), nuvärde:  
125 000 valutaenheter.  
Vilket räntebelopp ska du betala det andra året (d.v.s. i perioderna 13 till 24)?  
=KUMRÄNTA_ADD( 0,0075;360;125000;13;24;0) returnerar -11135,23.  
Hur mycket ränta måste du betala den första månaden?  
=KUMRÄNTA_ADD( 0,0075;360;125000;1;1;0) returnerar -937,50  
PRIS  
Beräknar värdet på ett värdepapper med fast ränta och det nominella värdet 100 valutaenheter oberoende av den avsedda avkastningen.  
Syntax  
PRIS( Betalning;Förfallodag;Ränta;Avkastning; Inlösningsvärde;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Ränta: den årliga nominella räntan (kupongränta).  
Avkastning: den årliga avkastningen på värdepapperet.  
Inlösningsvärde: inlösningsvärdet per 100 valutaenheter nominellt värde.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 15 februari 1999; förfallodagen är den 15 november 2007.  
Den nominella räntan är 5,75%.  
Avkastningen uppgår till 6,5%.  
Inlösningsvärdet ligger på 100 valutaenheter.  
Räntorna betalas halvårsvis (Frekvens är 2).  
Priset är följande vid beräkning med bas 0:  
=PRIS( "1999-02-15"; "2007-11-15"; 0,0575; 0,065; 100; 2; 0) returnerar 95,04287.  
PRISDISK  
Beräknar priset per 100 valutaenheter nominellt värde för ett diskonterat värdepapper.  
Syntax  
PRISDISK( Betalning;Förfallodag;Diskonteringsränta;Inlösningsvärde;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Diskonteringsränta: diskontering av värdepapperet i procent.  
Inlösningsvärde: inlösningsvärdet per 100 valutaenheter nominellt värde.  
Exempel  
Ett värdepapper köps den 15 februari 1999; förfallodagen är den 1 mars 1999.  
Diskonteringsräntan är 5,75%.  
Inlösningsvärdet ligger på 100.  
Priset är följande vid beräkning med bas 2:  
=PRISDISK( "1999-02-15"; "1999-03-01"; 0,0525; 100; 2) returnerar 99,79583.  
PRISFÖRF  
Beräknar priset per 100 valutaenheter nominellt värde för ett värdepapper som ger räntor på förfallodagen.  
Syntax  
PRISFÖRF( Betalning;Förfallodag;Emission;Ränta;Avkastning; Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Emission: datum för värdepappersemissionen.  
Ränta: räntesatsen för värdepapperet på emissionsdagen.  
Avkastning: den årliga avkastningen på värdepapperet.  
Exempel  
Betalning:  
15 februari 1999, Förfallodag:  
13 april 1999, Emission:  
11 november 1998.  
Ränta:  
6,1 procent, Avkastning:  
6,1 procent, Bas:  
30 / 360 = 0.  
Priset beräknas på följande sätt:  
=PRISFÖRF( "1999-02-15" ;"1999-04-13" ;"1998-11-11"; 0,061; 0,061;0) returnerar 99,98449888.  
LÖPTID  
LÖPTID är en funktion inom finansmatematiken.  
Du beräknar antalet perioder för en investering så att ett bestämt värde erhålls.  
Syntax  
LÖPTID( RÄNTA; Nuvärde;Slutvärde)  
Ränta är en konstant.  
Räntesatsen beräknas på hela löptiden.  
Räntesatsen per period räknas ut genom division av räntesatsen med den beräknade löptiden.  
Du anger räntesatsen för en annuitet som räntesats / 12.  
Nuvärde är det nuvarande värdet (dagsvärdet).  
Nuvärdet utgörs av ett investerat belopp eller en naturaförmån av motsvarande värde.  
Du måste ange ett positivt belopp som värde på investeringen; det får inte vara 0 eller <0.  
Slutvärde är det förväntade värdet.  
Det anger alltså vilket värde investeringen förväntas få i framtiden.  
Exempel  
Vid en räntesats på 4,75%, ett nuvarande värde på 25 000 valutaenheter och ett framtida värde på 1 000 000 valutaenheter returneras en löptid på 79,49 betalningsperioder.  
Den periodiska betalningen räknas ut genom att det framtida värdet divideras med löptiden, alltså:  
1 000 000 / 79,49=12 580,20.  
RRI.  
LINAVSKR  
Beräknar den linjära avskrivningen av en tillgång över en period.  
Avskrivningen är densamma över hela avskrivningstiden.  
Syntax  
LINAVSKR( AV; RV; LL)  
AV är tillgångens anskaffningsvärde.  
RV är tillgångens restvärde vid livslängdens slut.  
LL är livslängden uttryckt i antalet avskrivningsperioder.  
Exempel  
En kontorsutrustning med ett anskaffningsvärde på 50 000 valutaenheter ska skrivas av årligen under 7 år.  
Restvärdet är uppskattat till 3 500 valutaenheter.  
LINAVSKR( 50000;3500;84) = 553,57 valutaenheter.  
Den periodiska månatliga avskrivningen av kontorsutrustningen uppgår till 553,57 valutaenheter.  
ÅRSAVSKR, DEGAVSKR, VDEGRAVSKR.  
MLÖPTID  
Beräknar den modifierade Macauley-löptiden för ett värdepapper i år.  
Syntax  
MLÖPTID( Betalning;Förfallodag;Nominell ränta;Avkastning;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Nominell ränta: den årliga nominella räntan (kupongränta).  
Avkastning: den årliga avkastningen på värdepapperet.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps 1 januari 2001; förfallodag är 1 januari 2006.  
Den nominella räntan är 8%.  
Avkastningen är 9,0%.  
Hur lång är den modifierade löptiden vid beräkning exakt på dagen (bas 3)?  
=MLÖPTID( "01-01-01"; "06-01-01"; 0,08; 0,09; 2; 3)  
NETNUVÄRDE  
Beräknar kapitalvärdet av en investering baserat på en diskonteringsfaktor vid periodisk betalning (nettonuvärdet).  
Syntax  
NETNUVÄRDE( ränta;värde 1;värde 2;...)  
ränta är diskonteringsfaktorn för en period.  
värde1;... är upp till 30 värden som representerar in - eller utbetalningar.  
Exempel  
Hur stort är nettonuvärdet av periodiska betalningar på respektive 345, 276 och -145 valutaenheter med en diskonteringsfaktor på 8,75%?  
NETNUVÄRDE( 8,75%;345;276;-145) = 437,87 valutaenheter.  
Nettonuvärdet uppgår till 437,87 valutaenheter.  
NUVÄRDE, IR, SLUTVÄRDE.  
NOMRÄNTA  
Beräknar de årliga nominella räntorna till en effektiv ränta.  
Syntax  
NOMRÄNTA( ER;P)  
ER är den effektiva räntan.  
P är antalet periodiska räntebetalningar per år.  
Exempel  
Hur stora är de årliga nominalräntorna vid en effektiv ränta på 13,5% och tolv ränteinbetalningar per år?  
NOMRÄNTA( 13,5%;12) = 12,73%.  
Den årliga nominalräntesatsen är 12,73%.  
EFFRÄNTA.  
NOMRÄNTA_ADD  
Beräknar den årliga nominella räntan baserat på den effektiva räntan och antalet räntebetalningar per år.  
Syntax  
NOMRÄNTA_ADD( Effektiv ränta;Perioder)  
Effektiv ränta: den årliga effektiva räntan.  
Perioder: antalet räntebetalningar per år.  
Exempel  
Vad uppgår den nominella räntan till vid 5,3543% effektiv ränta och betalning kvartalsvis?  
=NOMRÄNTA_ADD( 5,3543%; 4) returnerar 0,0525 eller 5,25%.  
BRÅK  
Omvandlar en notering, som har angivits som ett decimaltal, till ett tal uttryckt som ett bråk.  
Syntax  
BRÅK( Tal;Nämnare)  
Tal: ett decimaltal.  
Nämnare: heltal som används som nämnare i bråket.  
Exempel  
=BRÅK( 1,125;16) omvandlar till sextondelar.  
Detta returnerar 1,02 för 1 plus 2 / 16.  
=BRÅK( 1,125;8) omvandlar till åttondelar.  
Detta returnerar 1,1 för 1 plus 1 / 8.  
DECTAL  
Omvandlar en notering, som har angivits som ett bråk, till ett decimaltal.  
Syntax  
DECTAL( Tal;Nämnare)  
Tal: ett tal angivet som bråk.  
Nämnare: heltal som används som nämnare i bråket.  
Exempel  
=DECTAL( 1,02;16) står för 1 och 2 / 16.  
Detta returnerar 1,125.  
=DECTAL( 1,1;8) står för 1 och 1 / 8.  
Detta returnerar 1,125.  
MODIR  
Beräknar den modifierade internräntan för en investeringsserie.  
Syntax  
MODIR( värden; investering; återinvestering)  
Värden motsvarar matrisen eller cellreferensen till celler vars innehåll motsvarar betalningarna.  
Investering är räntesatsen för investeringarna (de negativa värdena i matrisen)  
Återinvestering är räntesatsen för återinvesteringen (de positiva värdena i matrisen)  
Exempel  
Vid ett cellinnehåll i cellerna A1=-5, A2=10, A3=15 och A4=8, liksom ett investeringsvärde på 0,5 och ett återinvesteringsvärde på 0,1 blir resultatet 94,16%.  
NOMAVK  
Beräknar avkastningen på ett värdepapper.  
Syntax  
NOMAVK( Betalning;Förfallodag;Ränta;Pris;Inlösningsvärde;Frekvens;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Ränta: den årliga räntesatsen.  
Pris: priset (köppriset) på värdepapperet per 100 valutaenheter nominellt värde.  
Inlösningsvärde: inlösningsvärdet per 100 valutaenheter nominellt värde.  
Frekvens: antalet räntebetalningar per år (1, 2 eller 4).  
Exempel  
Ett värdepapper köps den 15 december 1999.  
Det förfaller den 15 november 2007.  
Räntesatsen är 5,75%.  
Priset är 95,04287 valutaenheter per 100 enheter nominellt värde, inlösningsvärdet är 100 enheter.  
Hur hög är avkastningen?  
=NOMAVK( "1999-02-15"; "2007-11-15"; 0,0575 ;95,04287; 100; 2; 0) returnerar 0,065 eller 6,5 procent.  
NOMAVKDISK  
Beräknar den årliga avkastningen på ett diskonterat värdepapper.  
Syntax  
NOMAVKDISK( Betalning;Förfallodag; Pris;Inlösningsvärde;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Pris: priset (köppriset) på värdepapperet per 100 valutaenheter nominellt värde.  
Inlösningsvärde: inlösningsvärde per 100 valutaenheter nominellt värde.  
Exempel  
Ett diskonterat värdepapper köps den 15 februari 1999.  
Det förfaller den 1 mars 1999.  
Priset är 99,795 valutaenheter per 100 enheter nominellt värde, inlösningsvärdet är 100 enheter.  
Hur hög är avkastningen?  
=NOMAVKDISK( "1999-02-15"; "1999-03-01"; 99,795; 100; 2) returnerar 0,052823 eller 5,2823 procent.  
NOMAVKFÖRF  
Beräknar den årliga avkastningen på ett värdepapper vars räntor betalas på förfallodagen.  
Syntax  
NOMAVKFÖRF( Betalning;Förfallodag;Emission;Ränta;Pris;Bas)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Emission: datum för värdepappersemissionen.  
Ränta: räntesatsen för värdepapperet på emissionsdagen.  
Pris: priset (köppriset) på värdepapperet per 100 valutaenheter nominellt värde.  
Exempel  
Ett värdepapper köps den 15 mars 1999.  
Det förfaller den 3 november 1999.  
Emissionsdag var den 8 november 1998.  
Räntesatsen är 6,25%, priset ligger på 100,0123 enheter.  
Hur hög är avkastningen?  
=NOMAVKFÖRF( "1999-03-15"; "1999-11-03"; "1998-11-08"; 0,0625; 100,0123; 0) returnerar 0,060954 eller 6,0954 procent.  
BETALNING  
Beräknar de regelbundna betalningarna (annuiteter) för en investering vid konstant räntesats.  
Syntax  
BETALNING( ränta; Perioder; NUVÄRDE; Slutvärde; F)  
ränta är räntesatsen för en periods betalning.  
Perioder är betalningstiden angiven i antalet perioder.  
Nuvärde är det nuvarande värdet av varje betalning.  
Slutvärde (valfritt) är det slutliga värde (framtida värde) som ska uppnås när de periodiska betalningarna har avslutats.  
F (valfritt) fastställer den periodiska betalningens förfallotid.  
F=1 anger betalning i början och F=0 betalning i slutet av en period.  
Exempel  
Hur stor är den regelbundna betalningen vid en räntesats på 1,99% om betalningsperioden är 3 år och nuvärdet 25 000 valutaenheter?  
BETALNING( 1,99%;36;25000) = -979,25 valutaenheter.  
Det regelbundna månatliga beloppet är alltså 979,25 valutaenheter.  
NUVÄRDE, AMORT, RÄNTA, RBETALNING, SLUTVÄRDE, PERIODER.  
SSVXEKV  
Beräknar den årliga räntan av en statsskuldsväxel (Treasury Bill).  
En statsskuldsväxel köps på likviddagen och säljs på förfallodagen, som måste vara samma år, till det fulla nominella värdet.  
En diskonteringsränta dras av från köppriset.  
Syntax  
SSVXEKV( Betalning;Förfallodag;Diskonteringsränta)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Diskonteringsränta: den procentuella diskonteringsräntan vid köpet av värdepapperet.  
Exempel  
Betalning:  
31 mars 1999, Förfallodag:  
1 juni 1999, Diskonteringsränta:  
9,14 procent.  
Förräntningen för statsskuldsväxeln motsvarande ett värdepapper räknas ut på följande sätt:  
=SSVXEKV( "1999-03-31" ;"1999-06-01"; 0,0914) returnerar 0,094151 eller 9,4151 procent.  
SSVXPRIS  
Beräknar priset på en statsskuldsväxel (Treasury Bill) per 100 valutaenheter.  
Syntax  
SSVXPRIS( Betalning;Förfallodag; Diskonteringsränta)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Diskonteringsränta: den procentuella diskonteringsräntan vid köpet av värdepapperet.  
Exempel  
Betalning:  
31 mars 1999, Förfallodag:  
1 juni 1999, Diskonteringsränta:  
9 procent.  
Priset på statsskuldsväxeln beräknas på följande sätt:  
=SSVXPRIS( "1999-03-31" ;"1999-06-01"; 0,09) returnerar 98,45.  
SSVXRÄNTA  
Beräknar avkastningen på en statsskuldsväxel (Treasury Bill).  
Syntax  
SSVXRÄNTA( Betalning;Förfallodag;Pris)  
Betalning: datum för värdepappersköpet.  
Förfallodag: datum då värdepapperet förfaller.  
Pris: priset (köppriset) på statsskuldsväxeln per 100 valutaenheter nominellt värde.  
Exempel  
Betalning:  
31 mars 1999, Förfallodag:  
1 juni 1999, Pris:  
98,45 valutaenheter.  
Avkastningen på en statsskuldsväxel beräknas på följande sätt:  
=SSVXRÄNTA( "1999-03-31" ;"1999-06-01"; 98,45) returnerar 0,091417 eller 9,1417 procent.  
Till finansfunktionerna del 1  
Till finansfunktionerna del 3  
Parameter till funktionen DAGAR360  
Tolkningsbeteendet hos DAGAR360-funktionen ändrades i och med lanseringen av %PRODUCTNAME 5.2.  
Det innebär att om du gör en ny beräkning av dokument från tidigare versioner kan det uppstå andra resultat.  
I det här avsnittet betyder "Gammal:" beteendet hos äldre %PRODUCTNAME -versioner än 5.2 och "Ny: "beteendet fr.o.m. %PRODUCTNAME version 5.2.  
Information:  
Den sista dagen i månaden är, med undantag av februari, alltid den 30:e (den 31:e behandlas som den 30:e).  
Månaden februari behandlas speciellt.  
Förändringarna i detalj:  
Gammal: den tredje alternativa paramatern ej angiven, tolkades som ej lika med 0 (TRUE) (europeisk metod).  
Ny: den tredje alternativa paramatern inte angiven, tolkas nu som lika med 0 (FALSE) (US-metod (NASD)).  
Gammal: om det äldre datumet är den 28 / 2 under ett skottår, omvandlas det till den 29 / 2 om den tredje parametern anges och om den är FALSE.  
Ny: om det äldre datumet är den 28 / 2 under ett skottår, förblir det alltid den 28 / 2.  
Tabellen visar en sammanfattning.  
Datum  
Skottår  
Parameter 3Typ  
Gammal:  
Ny:  
28.2.  
ja  
FALSE  
blev till den 29:e  
förblir den 28:e  
28.2.  
nej  
FALSE  
blev till den 30:e  
blir till den 30:e  
29.2.  
ja  
FALSE  
blev till den 30:e  
blir till den 30:e  
28.2.  
ja  
TRUE  
förblev den 28:e  
förblir den 28:e  
28.2.  
nej  
TRUE  
förblev den 28:e  
förblir den 28:e  
29.2.  
ja  
TRUE  
förblev den 29:e  
förblir den 29:e  
Därutöver gäller följande:  
Om det yngre datumet är den 31:e och den tredje parametern är FALSE och det äldre datumet inte är den 30:e. (efter eventuell omvandling av den 28 / 2 / 29 / 2. eller 31:e), då sätts det yngre datumet räknemässigt till den 1:e i följande månad.  
Om det yngre datumet är den 31:e och den tredje parametern är TRUE eller det äldre datumet är den 30:e, då sätts det yngre datumet till den 30:e.  
Behandlingen är (Gammal: / Ny:) densamma, men på grund av det ändrade standardvärdet om den tredje parametern saknas kan resultatet ändras.  
Exempel  
Gammal: =DAGAR360( 00.03.01; 00.03.31) = 29  
Ny: =DAGAR360( 00.03.01; 00.03.31) = 30  
=DAGAR360( 00.03.01; 00.03.31; FALSE) = 30  
=DAGAR360( 00.03.01;00.03.31; TRUE) = 29  
=DAGAR360( 00.02.28;00.03.01) = 3  
Gammal: =DAGAR360( 28.02.00;01.03.00; FALSE) = 2  
Ny: =DAGAR360( 00.02.28;00.03.01; FALSE) = 3  
=DAGAR360( 00.02.28;00.03.01; TRUE) = 3  
Gammal: =DAGAR360( 00.02.29; 00.03.01) = 2  
Ny: =DAGAR360( 00.02.29; 00.03.01) = 1  
=DAGAR360( 00.02.29; 00.03.01; FALSE) = 1  
=DAGAR360( 00.02.29;00.03.01; TRUE) = 2  
Statistik: grupp 1  
SKÄRNINGSPUNKT  
Här kan Du beräkna regressionslinjens skärningspunkt med y-axeln.  
Syntax  
SKÄRNINGSPUNKT( data_y; data_x)  
data_y är gruppen med beroende mätvärden eller data.  
data_x är gruppen med oberoende mätvärden eller data.  
Använd namn, matriser eller referenser som innehåller tal.  
Du kan naturligtvis även ange tal direkt.  
Exempel  
För beräkning av skärningen används cellerna D3:D9 ur exempeltabellen som y-värden och cellerna C3:C9 ur exempeltabellen som x-värden.  
De inmatade värdena ser alltså ut på följande sätt:  
SKÄRNINGSPUNKT( D3:D9;C3:C9) = 2,15.  
Resultatet är alltså 2,15.  
RKV, PEARSON, REGR, EXPREGR, PREDIKTION, LUTNING, STDFELYX, TREND, EXPTREND  
ANTAL  
Här kan Du beräkna det antal tal som en argumentlista består av.  
När antalet bestäms tas ingen hänsyn till textinmatningar.  
De enskilda värdena adderas.  
Syntax  
ANTAL( värde 1; värde 2; ...värde 30)  
värde 1; värde 2,...värde 30 är de värden ur vilka antalet argument räknas fram.  
Exempel  
Posterna 2,4,6 och åtta i textfälten värde 1-4 ska räknas.  
ANTAL( 2;4;6;åtta) = 3.  
Antalet poster är alltså 3.  
ANTALV, DANTAL, DANTALV, MEDEL, SUMMA  
ANTALV  
Beräknar antalet tal som en argumentlista innehåller.  
När antalet bestäms tas hänsyn till textinmatningar.  
De enskilda värdena adderas.  
Någon hänsyn tas inte till tomma argument.  
Syntax  
ANTALV( värde 1; värde 2; ...värde 30)  
värde 1; värde 2,...värde 30 är de värden ur vilka antalet argument räknas fram.  
Exempel  
Posterna 2,4,6 och åtta i textfälten värde1-4 ska räknas.  
ANTALV( 2;4;6;åtta) = 4.  
Antalet poster är alltså 4.  
ANTAL, DANTAL, DANTALV, MEDEL, PRODUKT, SUMMA  
B  
Sannolikheten för ett försöksresultat med binominalfördelning beräknas.  
Syntax  
B( försök;sannolikhet;G_1;G_2)  
försök bestämmer antalet försök.  
sannolikhet bestämmer den enskilda sannolikheten för ett försöksresultat.  
G_1 bestämmer den nedre gränsen för antalet försök.  
G_2 (valfri) bestämmer den övre gränsen för antalet försök.  
Exempel  
Hur stor är sannolikheten att man vid 10 kast med en tärning får upp sexan exakt två gånger?  
Det ger följande formel:  
=B( 10; 1 / 6; 2) ger 29% sannolikhet.  
BINOMFÖRD  
RKV  
När du vill beräkna kvadraten på den Pearsonska korrelationskoefficienten anger du respektive värden i textfälten.  
Korrelationskoefficienten är ett mått på kvaliteten på den anpassning som en regression kan uppnå och kallas också determinationskoefficient.  
Syntax  
RKV( data_y; data_x)  
data_y.  
Datapunkter i en matris eller ett område.  
data_x.  
Datapunkter i en matris eller ett område.  
Exempel  
=RKV( A1:A20; B1:B20) beräknar determinationskoefficienten för de två dataposterna i kolumnerna A och B.  
SKÄRNINGSPUNKT, KORREL, KOVAR, PEARSON, REGR, EXPREGR, LUTNING, STDFELYX, TREND  
BETAINV  
Returnerar värden för en inverterad betafördelad slumpvariabel.  
Syntax  
BETAINV( tal;alfa;beta;start;slut)  
tal är det värde med vilken funktionen ska utvärderas över intervallet start till slut.  
alfa är en fördelningsparameter.  
beta är en fördelningsparameter.  
start (valfri) är den nedre avgränsningen för tal.  
slut (valfri) är den övre avgränsningen för tal.  
Exempel  
=BETAINV( 0,5; 5; 10) ger värdet 0,33.  
BETAFÖRD  
BETAFÖRD  
Beräknar sannolikhetsfördelningen för en betafördelad slumpvariabel.  
Syntax  
BETAFÖRD( tal;alfa;beta;start;slut)  
tal är det värde med vilken funktionen ska utvärderas över intervallet start till slut.  
alfa är en fördelningsparameter.  
beta är en fördelningsparameter.  
start (valfri) är den nedre avgränsningen för tal.  
slut (valfri) är den övre avgränsningen för tal.  
Exempel  
=BETAFÖRD( 0,75; 3; 4) ger värdet 0,96.  
BETAINV  
BINOMFÖRD  
Beräknar sannolikheterna ur en binominalfördelad slumpvariabel.  
Syntax  
BINOMFÖRD( x;försök;sannolikhet;K)  
x är antalet lyckade försök i försöksserie.  
försök är det totala antalet försök.  
sannolikhet är sannolikheten för att ett försök ska vara lyckat.  
K = 0 beräknar den enkla och K = 1 den kumulerade sannolikheten.  
Exempel  
=BINOMFÖRD( A1; 12; 0,5; 0) visar, om Du sätter in värdena 0 till 12 istället för A1, sannolikheten att Du ska få exakt det antal förekomster av krona som anges i A1 om Du kastar ett mynt 12 gånger.  
=BINOMFÖRD( A1; 12; 0,5; 1) visar för samma rad den kumulerade sannolikheten, dvs. för A1=4 sannolikheten för att krona ska förekomma 0, 1, 2, 3 eller 4 gånger (ej exkluderande Eller).  
B, FAKULTET, HYPGEOMFÖRD, KOMBIN, KRITBINOM, NEGBINOMFÖRD, PERMUT, SANNOLIKHET  
CHI2INV  
Beräknar för en viss fastställd signifikansnivå värdet för den därtill hörande (teoretiska) chi2-fördelningen, som inte får överskridas av den observerade fördelningen, om den provade hypotesen ska vara sann.  
Chi2-fördelningen är en fördelningsfunktion ur statistiken, som fungerar som utgångspunkt för det s k "chi2-testet".  
Vid detta test provas en hypotes:  
Om den betraktade slumpstorheten uppfyller den fastställda fördelningslagen (dvs chi2-fördelningen) är hypotesen uppfylld.  
Under förutsättningen att hypotesen är sann, bör alltså den observerade chi-kvadraten motsvara den hypotetiska och teoretiska chi2-fördelningen (åtminstone ungefär).  
Chi2 beräknas som summan av  
(observerat värde-väntevärde )^2 / väntevärde  
för alla värden.  
Eftersom chi2 är ett mått på den sanna (observerade) fördelningens avvikelse från den hypotetiska (teoretiska), avvisas hypotesen om det chi2-värde som räknats fram ur ett konkret stickprov överskrider ett visst kritiskt värde.  
Den finns också angiven i tabeller i matematiska uppslagsverk.  
Syntax  
CHI2INV( tal; frihetsgrader)  
tal är värdet på den signifikansnivå till vilken den kritiska storheten CHIINV ska beräknas, dvs den sannolikhet med vilken hypotesen är säkrad.  
frihetsgrader är antalet frihetsgrader i experimentet.  
Exempel  
En tärning kastas 1020 gånger.  
Antalet prickar, från 1 till 6, förekommer 195, 151, 148, 189, 183 respektive 154 gånger (observationsvärden).  
Det ska provas om tärningen är omanipulerad.  
Stickprovets chi2-fördelning beräknas med ovanstående formel.  
1020 / 6 = 170, ger formeln ett chi2-värde på 13,27.  
Om den (observerade) chi-kvadraten är större än eller lika med den (teoretiska) chi-kvadraten CH2INV, förkastas hypotesen, eftersom avvikelsen mellan teori och experiment är för stor.  
Om den observerade chi-kvadraten är mindre än CHI2INV godtas hypotesen med den angivna signifikansnivån.  
=CHI2INV( 0,05; 5) ger 11,07.  
=CHI2INV( 0,05; 5) ger 13,39.  
Med en signifikansnivå på 5% är tärningen inte omanipulerad, med en signifikansnivå på 2% finns det ingen orsak att betvivla att den skulle vara omanipulerad.  
CHI2TEST, CHI2FÖRD  
CHI2TEST  
Ger med hjälp av chi2-testet ur mätdata direkt sannolikhetsvärdet för att en hypotes är uppfylld.  
Observerade och förväntade storheter i ett stickprov jämförs:  
CHI2TEST jämför de båda dataraderna och beräknar Chi2-värdet ur summan av (observerat värde-förväntat värde )^2 / förväntat värde för alla värden.  
Ur detta chi2-värde beräknas slutligen signifikansnivån hos den hypotes som ska provas.  
Istället för datakolumnerna ska stickprovets chi-kvadrat överlämnas som parameter.  
Syntax  
CHI2TEST( data_B; data_F)  
data_B är matrisen med de observerade värdena.  
data_F är matrisen med de förväntade värdena.  
Exempel  
A (observerad)  
B (förväntad)  
1  
195  
170  
2  
151  
170  
3  
148  
170  
4  
189  
170  
5  
183  
170  
6  
154  
170  
=CHI2TEST( A1:A6; B1:B6) ger 0,02.  
Det är sannolikheten med vilka observerade data uppfyller den teoretiska chi2-fördelningen.  
CHI2INV, CHI2FÖRD  
CHI2FÖRD  
Ger ur den angivna chi-kvadraten sannolikhetsvärdet för att en hypotes är uppfylld.  
Ur detta fastställs signifikansnivån för den provade hypotesen.  
Istället för stickprovets chi-kvadrat ska observerade och förväntade data överlämnas som parametrar.  
Syntax  
CHI2FÖRD( tal; frihetsgrader)  
tal är stickprovets chi2-värde, till vilken signifikansnivån ska beräknas.  
frihetsgrader är antalet frihetsgrader i experimentet.  
Exempel  
=CHI2FÖRD( 13,27; 5) ger 0,02.  
Om stickprovets chi2-värde uppgår till 13,27 och om experimentet har 5 frihetsgrader är hypotesen säkerställd med en signifikansnivå på 2%.  
CHI2INV, CHI2TEST  
EXPONFÖRD  
Beräknar sannolikheten för en exponentialfördelad slumpvariabel.  
Syntax  
EXPONFÖRD( tal; lambda; kumulativ)  
tal är det värde för vilket exponentialfördelningen ska beräknas.  
lambda är exponentialfördelningens parameter.  
kumulativ K = 0 beräknar täthetsfunktionen, K = 1 fördelningen.  
Exempel  
=EXPONFÖRD( 3; 0,5; 1) ger 0,78.  
GAMMAFÖRD, POISSON  
Statistik: grupp 2  
FINV  
Beräknar inversen på F-fördelningen.  
F-fördelningen används i F-tester för att bestämma sambandet mellan två datamängder med var sin fördelning.  
Syntax  
FINV( tal; frihetsgrader_1; frihetsgrader_2)  
tal är sannolikhetsvärdet för vilket den inverterade F-fördelningen ska beräknas.  
frihetsgrader_1 är antalet frihetsgrader i F-fördelningens täljare.  
frihetsgrader_2 är antalet frihetsgrader i F-fördelningens nämnare.  
Exempel  
=FINV( 0,5; 5; 10) ger 0,93.  
FTEST, FFÃ–RD  
FISHER  
Räknar igenom Fisher-transformationen för x och skapar en funktion som är ganska normalfördelad och därmed besitter en snedhet på ungefär 0.  
Syntax  
FISHER( tal)  
tal är värdet som ska transformeras.  
Exempel  
=FISHER( 0,5) ger 0,55.  
FISHERINV, KORREL, KOVAR  
FISHERINV  
Räknar igenom Fisher-transformationen inverterat för x och skapar en funktion som är ganska normalfördelad och därmed besitter en snedhet på ungefär 0.  
Syntax  
FISHERINV( tal)  
tal är värdet som ska återtransformeras.  
Exempel  
=FISHERINV( 0,5) ger 0,46.  
FISHER, KORREL, KOVAR  
FTEST  
Genomför en F-varianstest och beräknar statistiken.  
Syntax  
FTEST( data_1; data_2)  
data_1 är den första datapostens matris.  
data_2 är den andra datapostens matris.  
Exempel  
=FTEST( A1:A30; B1:B12) beräknar om de två datakolumnerna skiljer sig åt i varians och ger som resultat hur sannolikt det är att de två kolumnerna kommer från samma population.  
FINV, FFÃ–RD  
FFÖRD  
Beräknar F-fördelningsfunktionens värden.  
Syntax  
FFÖRD( tal; frihetsgrader_1; frihetsgrader_2)  
tal är värdet för vilket F-fördelningen ska beräknas.  
frihetsgrader_1 är antalet frihetsgrader i F-fördelningens täljare.  
frihetsgrader_2 är antalet frihetsgrader i F-fördelningens nämnare.  
Exempel  
=FFÖRD( 0,8; 8; 12) ger 0,61.  
FINV, FTEST  
GAMMAINV  
Beräknar inversen på gammafördelningen.  
Med denna funktion kan Du undersöka variabler vars fördelning eventuellt är ojämna.  
Syntax  
GAMMAINV( tal; alfa; beta)  
tal är sannolikhetsvärdet för vilket den inversa gammafördelningen ska beräknas.  
alfa är gammafördelningens alfaparameter.  
beta är gammafördelningens betaparameter.  
Exempel  
=GAMMAINV( 0,8; 1; 1) ger 1,61.  
GAMMAFÖRD  
GAMMALN  
Beräknar Gamma-funktionens naturliga logaritm G( x).  
Syntax  
GAMMALN( tal)  
tal är värdet för vilket Gamma-funktionens naturliga logaritm ska beräknas.  
Exempel  
=GAMMALN( 2) ger 0.  
FAKULTET  
GAMMAFÖRD  
Beräknar sannolikheten för en gammafördelad slumpvariabel.  
Syntax  
GAMMAFÖRD( tal; alfa; beta; kumulativ)  
tal är värdet för vilket gammafördelningen ska beräknas.  
alfa är gammafördelningens alfaparameter.  
beta är gammafördelningens alfaparameter.  
kumulativ = 0 beräknar täthetsfunktionen, kumulativ = 1 fördelningen.  
Exempel  
=GAMMAFÖRD( 0,8; 1; 1) ger 0,86.  
CHI2FÖRD, EXPONFÖRD, GAMMAINV  
GAUSS  
Bestämmer standardnormalfördelningens integralvärde.  
Syntax  
GAUSS( tal)  
tal är värdet för vilket standardnormalfördelningens integralvärde ska beräknas.  
Exempel  
GAUSS( 0,19) = 0,08  
GAUSS( 0,0375) = 0,01  
ZTEST, NORMFÖRD, NORMSFÃ–RD  
GEOMEAN  
Beräknar det geometriska medelvärdet för en mängd positiva tal.  
Syntax  
GEOMEAN( tal 1; tal 2; ...tal 30)  
tal 1, tal 2,...tal 30 är numeriska argument som representerar ett stickprov.  
Exempel  
Om Du skriver in värdena 23, 46 och 69 i textfälten tal 1, 2 och 3 får Du 41,79 som resultat.  
GEOMEAN( 23; 46; 69) = 41,79.  
Det här stickprovets geometriska medelvärde är alltså 41,79.  
TRIMMEDEL, HARMMEDEL, MEDIAN, MEDEL, TYPVÄRDE  
TRIMMEDEL  
Beräknar en datagrupps medelvärde, utan att ta hänsyn till värdena vid kanterna.  
Syntax  
TRIMMEDEL( data; alfa)  
data är datamatrisen i stickprovet.  
alfa är procentsatsen för marginalvärdena som det inte ska tas någon hänsyn till.  
Exempel  
=TRIMMEDEL( A1:A50;0,1) beräknar medelvärdet för talen i A1:A50, utan att ta hänsyn till de 5% lägsta och de 5% högsta värdena.  
Procenttalen hänför sig till värdet för det otrimmade medelvärdet och inte antalet summander.  
GEOMEAN, HARMMEDEL, MEDIAN, MEDEL, TYPVÄRDE  
ZTEST  
Beräknar den tvåsidiga kontrollstatistiken för ett Gausstest med normalfördelning.  
Syntax  
ZTEST( data; x; STD)  
data är datamatrisen.  
x är det värde som ska testas.  
STD (valfri) är populationens standardavvikelse.  
Saknas detta argument görs beräkningarna med respektive stickprovs standardavvikelse.  
Exempel  
=ZTEST( A1:A50; 12) ger sannolikheten för att värdet 12 hör till den normalfördelade populationen i A1:A50.  
KONFIDENS, NORMINV, NORMFÖRD, STANDARDISERA, NORMSINV, NORMSFÖRD  
HARMMEDEL  
Beräknar en datamängds harmoniska medelvärde.  
Syntax  
HARMMEDEL( tal 1; tal 2; ...tal 30)  
tal 1,tal 2,...tal 30 är upp till 30 argument som används för att beräkna det harmoniska medelvärdet.  
Exempel  
Om Du matar in värdena 23, 46 och 69 i textfälten tal 1, 2 och 3 får Du 37,64 som resultat.  
HARMMEDEL( 23;46;69) = 37,64.  
Det harmoniska medelvärdet för detta stickprov är alltså 37,64.  
GEOMEAN, TRIMMEDEL, MEDIAN, MEDEL, TYPVÄRDE  
HYPGEOMFÖRD  
Beräknar sannolikheten i hypergeometriskt fördelade slumpvariabler.  
Syntax  
HYPGEOMFÖRD( X; storlek; population; populationsstorlek)  
X är antalet lyckade försök i stickprovet.  
storlek är stickprovets storlek.  
population är antalet lyckade försök i populationen.  
populationsstorlek är populationens storlek.  
Exempel  
=HYPGEOMFÖRD( 2; 2; 90; 100) ger 0,81.  
Om 90 av 100 smörgåsar ramlar med smörsidan nedåt från bordet och om jag låter två smörgåsar falla från bordet, är sannolikheten 81% för att båda smörgåsarna ska hamna med smörsidan nedåt.  
BINOMFÖRD, FAKULTET, KOMBIN, NEGBINOMFÖRD, PERMUT  
Statistik: grupp 3  
STÖRSTA  
Beräknar det k:te största värdet i en datagrupp.  
Syntax  
STÖRSTA( data; rang_k)  
data är datamatrisen i stickprovet.  
rang_k är värdets rangordning.  
Exempel  
=STÖRSTA( A1:C50; 2) ger det näst största värdet i A1:C50.  
MINSTA, MAX, MEDIAN, PERCENTIL, PROCENTRANG, KVARTIL  
MINSTA  
Beräknar det k:te minsta värdet i en datagrupp.  
Syntax  
MINSTA( data; rang_k)  
data är datamatrisen i stickprovet.  
rang_k är värdets rangordning.  
Exempel  
=MINSTA( A1:C50; 2) ger det näst minsta värdet i A1:C50.  
STÖRSTA, MEDIAN, MIN, PERCENTIL, PROCENTRANG, KVARTIL  
KONFIDENS  
Beräknar ett (1-alfa) konfidensintervall för normalfördelningen.  
Syntax  
KONFIDENS( alfa; STD; storlek)  
alfa är konfidensintervallets nivå.  
STD är populationens standardavvikelse.  
N är populationens storlek.  
Exempel  
=KONFIDENS( 0,05; 1,5; 100) ger 0,29.  
ZTEST  
KORREL  
Beräknar en tvådimensionell slumpstorhets korrelationskoefficient.  
Syntax  
KORREL( data_1; data_2)  
data_1 är den första datapostens matris.  
data_2 är den andra datapostens matris.  
Exempel  
=KORREL( A1:A50; B1:B50) beräknar korrelationskoefficienten som ett mått på det linjära sambandet mellan de två datakolumnerna.  
FISHER, FISHERINV, KOVAR  
KOVAR  
Beräknar kovariansen för alla produkter som bildats i datapunktsparen.  
Syntax  
KOVAR( data_1; data_2)  
data_1 är den första datapostens matris.  
data_2 är den andra datapostens matris.  
Exempel  
=KOVAR( A1:A30; B1:B30)  
FISHER, FISHERINV, KORREL  
KRITBINOM  
Beräknar det minsta värde för vilket den kumulerade sannolikheten hos binominalfördelningen är lika med eller större än en viss gränssannolikhet.  
Syntax  
KRITBINOM( försök; sannolikhet; alfa)  
försök är det totala antalet försök.  
sannolikhet är sannolikheten för att ett försök ska vara lyckat.  
alfa är gränssannolikheten som ska uppnås eller överskridas.  
Exempel  
=KRITBINOM( 100; 0,5; 0,1) ger 44.  
BINOMFÖRD, FAKULTET, HYPGEOMFÖRD, KOMBIN, NEGBINOMFÖRD, PERMUT, SANNOLIKHET  
TOPPIGHET  
Beräknar en datagrupps kurtosis (excess).  
Du måste skriva in minst 4 värden.  
Syntax  
TOPPIGHET( tal 1; tal 2; ...tal 30)  
tal 1, tal 2,...tal 30 är numeriska argument som representerar ett stickprov i fördelningen.  
Exempel  
=TOPPIGHET( A1;A2;A3;A4;A5;A6)  
SNEDHET, STDAV, STDAVP, VARIANS, VARIANSP  
LOGINV  
Beräknar den logaritmiska normalfördelningens inverterade funktion.  
Syntax  
LOGINV( tal; MV; STD)  
tal är sannolikhetsvärdet för vilket den inversa lognormalfördelningen ska beräknas.  
MV är lognormalfördelningens medelvärde.  
STD är standardavvikelsen från lognormalfördelningen.  
Exempel  
=LOGINV( 0,05; 0; 1) ger 0,19.  
EXP, LN, LOG, LOG10, LOGNORMFÃ–RD  
LOGNORMFÖRD  
Beräknar fördelningsfunktionens värden hos en lognormfördelad slumpvariabel.  
Syntax  
LOGNORMFÖRD( tal; MV; STD)  
tal är sannolikhetsvärdet för vilket lognormalfördelningen ska beräknas.  
MV är lognormalfördelningens medelvärde.  
STD är standardavvikelsen från lognormalfördelningen.  
Exempel  
=LOGNORMFÖRD( 0,1; 0; 1) ger 0,01.  
EXP, LN, LOG, LOG10, LOGINV  
Statistik: grupp 4  
MAX  
Beräknar det största värdet inom en argumentlista.  
Syntax  
MAX( tal 1; tal 2; ...tal 30)  
tal 1; tal 2 ;...tal 30 är numeriska argument, vars största tal ska bestämmas.  
Vart och ett av talen kan även ersättas med en referens.  
Exempel  
=MAX( A1;A2;A3;50;100;200) returnerar det största värdet från den här listan.  
=MAX( A1:B100) returnerar det största värdet från den här listan.  
DMAX, MIN  
MAXA  
Beräknar det största värdet inom en argumentlista.  
Texten värderas då till 0.  
Syntax  
MAXA( värde 1; värde 2; ...värde 30)  
värde 1; värde 2 ;...värde 30 är de argument, vars största värde ska bestämmas.  
Vart och ett av värdena kan även ersättas med en referens.  
En text värderas då som 0.  
Exempel  
=MAXA( A1;A2;A3;50;100;200) returnerar det största värdet från den här listan.  
=MAXA( A1:B100) returnerar det största värdet från den här listan.  
MINA  
MEDIAN  
Beräkna medianen (mittpunkten) för de angivna talen.  
För en talserie med ojämnt antal är medianen det värde som står mitt i listan.  
För en talserie med jämnt antal beräknas medelvärdet för det två mellersta värdena.  
Syntax  
MEDIAN( tal 1; tal 2; ...tal 30)  
tal 1; tal 2 ;...tal 30 är argument, som utgör ett stickprov.  
Vart och ett av talen kan även ersättas med en referens.  
Exempel  
(udda antal): =MEDIAN(1, 5, 9, 20, 21) returnerar det mellersta värdet från den här listan, d v s 9.  
(jämnt antal): =MEDIAN(1, 5, 9, 20) returnerar medelvärdet för de båda mellersta värdena 5 och 9, d v s 7.  
ANTAL, ANTALV, DMEDEL, MEDEL, TYPVÄRDE, SUMMA  
MIN  
Returnerar det minsta talet i en lista med argument.  
Syntax  
MIN( tal 1; tal 2; ...tal 30)  
tal 1; tal 2 ;...tal 30 är numeriska argument, vars minsta tal ska bestämmas.  
Vart och ett av talen kan även ersättas med en referens.  
Exempel  
=MIN( A1:B100) returnerar det minsta värdet från den här listan.  
DMIN, MAX  
MINA  
Returnerar det minsta värdet från en lista med argument.  
Förutom tal kan även text anges.  
Text värderas till 0.  
Syntax  
MINA( värde 1; värde 2; ...värde 30)  
värde 1; värde 2 ;...värde 30 är de argument, vars minsta värde ska bestämmas.  
Vart och ett av värdena kan även ersättas med en referens.  
Text värderas till 0.  
Exempel  
=MINA( 1; text; 20) returnerar det minsta värdet från den här listan.  
=MINA( A1:B100) returnerar det minsta värdet från den här listan.  
MAXA  
MEDELAVV  
Returnerar medelvärdet för datapunkters absoluta avvikelse från deras medelvärde.  
Visar spridningen i ett dataområde.  
Syntax  
MEDELAVV( tal 1; tal 2; ...tal 30)  
tal 1; tal 2 ;...tal 30 är argument, som utgör ett stickprov.  
Vart och ett av talen kan även ersättas med en referens.  
Exempel  
=MEDELAVV( A1:A50)  
STDAV, STDAVP, KVADAVV, VARIANS, VARIANSP  
MEDEL  
Beräknar det aritmetiska medelvärdet för argumenten.  
Syntax  
MEDEL( tal 1; tal 2; ...tal 30)  
tal 1; tal 2 ;...tal 30 är numeriska argument som utgör ett stickprov taget ur en population.  
Vart och ett av talen kan även ersättas med en referens.  
Exempel  
=MEDEL( A1:A50)  
GEOMEDEL, TRIMMEDEL, HARMMEDEL, MEDIAN, TYPVÄRDE  
MEDELA  
Beräknar det aritmetiska medelvärdet för argumenten.  
Text värderas till 0.  
Syntax  
MEDELA( värde 1; värde 2; ...värde 30)  
värde 1; värde 2 ;...värde 30 är argument som utgör ett stickprov taget ur en population.  
Vart och ett av värdena kan även ersättas med en referens.  
Text värderas till 0.  
Exempel  
=MEDELA( A1:A50)  
MEDEL  
TYPVÄRDE  
Returnerar det värde som oftast förekommer i en matris eller i ett dataområde.  
Om det finns flera värden med samma frekvens returneras det minsta av dessa.  
Om inget värde förekommer två gånger returneras ett felmeddelande.  
Syntax  
TYPVÄRDE( tal 1; tal 2; ...tal 30)  
tal 1; tal 2 ;...tal 30 är numeriska argument som utgör ett stickprov.  
Vart och ett av talen kan även ersättas med en referens.  
Exempel  
=TYPVÄRDE( A1:A50)  
GEOMEDEL, TRIMMEDEL, HARMMEDEL, MEDIAN, MEDEL  
NEGBINOMFÖRD  
Returnerar sannolikheten för en negativt binomialfördelad slumpvariabel.  
Syntax  
NEGBINOMFÖRD( x; R; sannolikhet)  
x är antalet misslyckanden i försöksserien.  
R är antalet lyckade försök i serien.  
sannolikhet är sannolikheten för ett lyckat försök.  
Exempel  
=NEGBINOMFÖRD( 1; 1; 0,5) ger resultatet 0,25.  
BINOMFÖRD, FAKULTET, HYPGEOMFÖRD, KOMBIN, PERMUT  
NORMINV  
Returnerar normalfördelningens del för det angivna medelvärdet och standardavvikelsen.  
Syntax  
NORMINV( tal; MV; STD)  
tal är sannolikhetsvärdet för vilket den inversa normalfördelningen ska beräknas.  
MV är medelvärdet för normalfördelningen.  
STD är standardavvikelsen för normalfördelningen.  
Exempel  
=NORMINV( 0,9; 63; 5) ger resultatet 69,41.  
Om ett standardfrukostägg väger 63 g, med en standardavvikelse på 5, så väger ägget med 90% sannolikhet max 69,41 g.  
ZTEST, NORMFÖRD, STANDARDISERA, NORMSINV, NORMSFÖRD  
NORMFÖRD  
Returnerar sannolikheterna för en normalfördelad slumpvariabel för det angivna medelvärdet och standardavvikelsen.  
Syntax  
NORMFÖRD( tal; MV; STD; K)  
tal är det fördelningsvärde för vilket normalfördelningen ska beräknas.  
MV är det aritmetiska medelvärdet för fördelningen.  
STD är standardavvikelsen för fördelningen.  
K = 0 returnerar frekvensfunktionen, K = 1 returnerar fördelningen.  
Exempel  
=NORMFÖRD( 70; 63; 5; 0) ger resultatet 0,03.  
=NORMFÖRD( 70; 63; 5; 1) ger resultatet 0,92.  
ZTEST, NORMINV, STANDARDISERA, NORMSINV, NORMSFÖRD  
PEARSON  
Returnerar Pearsons korrelationskoefficient r.  
Syntax  
PEARSON( data_1; data_2)  
data_1 är den första datapostens matris.  
data_2 är den andra datapostens matris.  
Exempel  
=PEARSON( A1:A30; B1:B30) returnerar Pearsons korrelationskoefficient för de båda dataserierna.  
SKÄRNINGSPUNKT, RKV, REGR, LUTNING, STDFELYX  
PHI  
Returnerar värdet av fördelningsfunktionen för standardnormalfördelningen.  
Syntax  
PHI( tal)  
tal är värdet för vilket standardnormalfördelningen beräknas.  
Exempel  
PHI( 2,25) = 0,03  
PHI( -2,25) = 0,03  
PHI( 0) = 0,4  
NORMSFÖRD  
POISSON  
Beräkna sannolikheten för en Poisson-fördelad slumpvariabel.  
Syntax  
POISSON( tal; MV; K)  
tal är värdet för vilket Poisson-fördelningen ska beräknas.  
MV är medelvärdet för Poisson-fördelningen.  
K = 0 returnerar frekvensfunktionen, K = 1 returnerar fördelningen.  
Exempel  
=POISSON( 60;50;1) ger resultatet 0,93.  
EXPONFÖRD  
PERCENTIL  
Beräknar en alfa-kvantil för ett stickprov.  
En percentil returnerar ett skalvärde för en dataserie, som ligger på alfa procent av skalan från det minsta till det största värdet i dataserien.  
För alfa = 25% kallas percentilen första kvartilen, för alfa = 50% kallas den MEDIAN.  
Syntax  
PERCENTIL( data;alfa)  
data är datamatrisen.  
alfa definierar procentsatsen för percentilen, som ligger mellan 0 och 1.  
Exempel  
=PERCENTIL( A1:A50; 0,1) returnerar det värde i dataserien, som utgör 10% av totala spannet för alla data inom A1:A50:  
STÖRSTA, MINSTA, MAX, MEDIAN, MIN, PROCENTRANG, KVARTIL  
PROCENTRANG  
Beräknar den procentuella rangen (alfa) för ett värdet i ett stickprov.  
Syntax  
PROCENTRANG( data; värde)  
data är datamatrisen i stickprovet.  
värde är det värde, vars procentuella rang ska bestämmas.  
Exempel  
=PROCENTRANG( A1:A50; 50) returnerar den procentuella rangen för värdet 50 i det totala området för alla värden inom A1:A50.  
Om 50 ligger utanför det totala området visas ett felmeddelande.  
STÖRSTA, MINSTA, MAX, MEDIAN, MIN, PERCENTIL, KVARTIL  
KVARTIL  
Beräknar kvartilen för ett stickprov.  
Syntax  
KVARTIL( data; typ)  
data är datamatrisen i stickprovet.  
typ är typen av kvartil. (0 = MIN, 1 = 25%, 2 = 50% (MEDIAN), 3 = 75% och 4 = MAX.)  
Exempel  
=KVARTIL( A1:A50; 2) returnerar det värde som motsvarar 25% av skalan från minsta till största värdet i området A1:A50.  
STÖRSTA, MINSTA, MAX, MEDIAN, MIN, PERCENTIL, PROCENTRANG  
Statistik: grupp 5  
RANG  
Beräknar rangen för ett värde i ett stickprov.  
Syntax  
RANG( värde; data; typ)  
värde är värdet vars rang ska bestämmas.  
data är datamatrisen i stickprovet.  
typ (valfri) är ordningsföljden som används i rangordningen. typ=0 betyder stigande, typ=1 betyder fallande.  
Exempel  
=RANG( A10; A1:A50) ger rangplaceringen för värdet i A10 inom värdena i området A1:A50.  
Om värde inte finns i området visas ett felmeddelande.  
PROCENTRANG  
SNEDHET  
Beräknar den matematiska snedheten för en fördelning.  
Syntax  
SNEDHET( tal 1; tal 2; ...tal 30)  
tal 1, tal 2...tal 30 är numeriska argument som utgör stickprov för fördelningen.  
Du kan även ange områden.  
Exempel  
=SNEDHET( A1:A50) beräknar värdet på snedheten för data i den angivna referensen.  
TOPPIGHET, STDAV, STDAVP, VARIANS, VARIANSP  
PREDIKTION  
Beräknar ett värde längs en regressionslinje.  
Syntax  
PREDIKTION( värde; data_y; data_x)  
värde är x-värdet för vilket y-värdet på regressionslinjen ska beräknas.  
data_y är matrisen med y-data.  
data_x är matrisen med x-data.  
Exempel  
=PREDIKTION( 50; A1:A50; B1;B50) returnerar det y-värde som förväntas för x-värdet 50 om x - och y-värdena i de båda referenserna är kopplade med linjär regression.  
REGR, EXPREGR, TREND, EXPTREND  
STDAV  
Beräknar standardavvikelsen baserad på ett stickprov.  
Syntax  
STDAV( tal 1;tal 2;...tal 30)  
tal 1, tal 2...tal 30 är numeriska argument som utgör ett stickprov från en population.  
Exempel  
=STDAV( A1:A50) returnerar den uppskattade standardavvikelsen baserad på data i referensen.  
MEDELAVV, MEDEL, TYPVÄRDE, STDAVP, VARIANS  
STDAVA  
Beräknar standardavvikelsen baserat på ett stickprov.  
Text värderas till 0.  
Syntax  
STDAVA( värde 1;värde 2;...värde 30)  
värde 1, värde 2...värde 30 är argument som utgör ett stickprov ur en population.  
Texter är också möjliga och värderas till 0.  
Exempel  
=STDAVA( A1:A50) returnerar den uppskattade standardavvikelsen baserat på data i referensen.  
STDAV, STDAVP och STDAVPA.  
STDAVP  
Beräknar standardavvikelsen baserat på populationen.  
Syntax  
STDAVP( tal 1;tal 2;...tal 30)  
tal 1, tal 2...tal 30 är numeriska argument som utgör ett stickprov från en population.  
Exempel  
=STDAVP( A1:A50) returnerar standardavvikelsen baserat på data i referensen.  
MEDELAVV, MEDEL, TYPVÄRDE, STDAV, VARIANSP  
STDAVPA  
Beräknar standardavvikelsen baserat på populationen.  
Text värderas till 0.  
Syntax  
STDAVPA( värde 1;värde 2;...värde 30)  
värde 1, värde 2...värde 30 är argument som utgör stickprov ur en population.  
Text värderas till 0.  
Exempel  
=STDAVPA( A1:A50) returnerar standardavvikelsen baserad på data i referensen.  
STDAVP och STDAVA.  
STANDARDISERA  
Beräknar det standardiserade värdet för en fördelning kännetecknad av medelvärde och standardavvikelse.  
Syntax  
STANDARDISERA( tal; MV; STD)  
tal är värdet som ska standardiseras.  
MV är medelvärdet med vilket förflyttningen ska göras.  
STD är standardavvikelsen med vilket skalningen ska göras.  
Exempel  
=STANDARDISERA( 11; 10; 1) returnerar 1.  
Värdet 11 ligger i en normalfördelning med medelvärdet 10 och standardavvikelsen 1 lika långt över medelvärdet 10 som värdet 1 ligger över medelvärdet 0 i standardnormalfördelningen.  
ZTEST, NORMINV, NORMFÖRD, NORMSINV, NORMSFÖRD  
NORMSINV  
Beräknar värden för den inversa standardnormalfördelningen.  
Syntax  
NORMSINV( tal)  
tal är sannolikhetsvärdet för vilket den inversa standardnormalfördelningen ska beräknas.  
Exempel  
NORMSINV( 0,908789) returnerar 1,3333.  
ZTEST, NORMINV, NORMFÖRD, STANDARDISERA, NORMSFÖRD  
NORMSFÖRD  
Beräknar värdet av fördelningsfunktionen för standardnormalfördelade slumpvariabler.  
Syntax  
NORMSFÖRD( tal)  
tal är det värde för vilket standardnormalfördelningen ska beräknas.  
Exempel  
=NORMSFÖRD( 1) returnerar 0,84.  
Det betyder att ytan under standardnormalfördelningens kurva till vänster om x-värdet 1 utgör 84% av den totala ytan.  
ZTEST, NORMINV, NORMFÖRD, PHI, STANDARDISERA, NORMSINV  
LUTNING  
Beräknar lutningen på en linjär regressionslinje.  
Den anpassas till de datapunkter som har lagrats i x - och y-värdena.  
Syntax  
LUTNING( data_y; data_x)  
data_y är matrisen med y-data.  
data_x är matrisen med x-data.  
Exempel  
=LUTNING( A1:A50; B1:B50)  
SKÄRNINGSPUNKT, RKV, PEARSON, REGR, EXPREGR, STDFELYX, TREND  
STDFELYX  
Beräknar standardfelet i de uppskattade y-värdena för varje x-värde i regressionen.  
Syntax  
STDFELYX( data_y; data_x)  
data_y är matrisen med y-data.  
data_x är matrisen med x-data.  
Exempel  
=STDFELXY( A1:A50; B1:B50)  
SKÄRNINGSPUNKT, RKV, PEARSON, REGR, EXPREGR, LUTNING  
KVADAVV  
Beräknar summan av den kvadratiska avvikelsen hos datapunkter från ett stickprovs medelvärde.  
Syntax  
KVADAVV( tal 1; tal 2; ...tal 30)  
tal 1, tal 2...tal 30 är numeriska argument som utgör ett stickprov.  
Du kan även ange referenser.  
Exempel  
=KVADAVV( A1:A50)  
MEDELAVV, STDAV, STDAVP, VARIANS, VARIANSP  
TINV  
Beräknar värden för den inversa (Students) t-fördelningen för de angivna frihetsgraderna.  
Syntax  
TINV( tal; frihetsgrader)  
tal är sannolikhetsvärdet för vilket den inversa t-fördelningen ska beräknas.  
frihetsgrader är antalet frihetsgrader i t-fördelningen.  
Exempel  
=TINV( 0,1; 6) returnerar 1,94  
TTEST, TFÖRD  
TTEST  
Beräknar teststatistiken för en students t-test.  
Syntax  
TTEST( data_1; data_2; läge; typ)  
data_1 är matrisen för den första dataposten.  
data_2 är matrisen för den andra dataposten.  
läge = 1 beräknar det ensidiga testet, läge = 2 det tvåsidiga.  
Typ 1 betyder parad.  
Typ 3 betyder två stickprov med olika varians (heteroskedastisk).  
Exempel  
=TTEST( A1:A50; B1:B50; 2; 2)  
TINV, TFÖRD  
TFÖRD  
Beräknar värdet på fördelningsfunktionen (1-alfa) för en (students) t-fördelade slumpvariabel.  
Syntax  
TFÖRD( tal; frihetsgrader; läge)  
tal är det värde för vilket t-fördelningen ska beräknas.  
frihetsgrader är frihetsgraderna i t-fördelningen.  
läge = 1 beräknar det ensidiga testet, läge = 2 det tvåsidiga.  
Exempel  
=TFÖRD( 12; 5; 1)  
TINV, TTEST  
Varians  
Beräknar en uppskattning av variansen baserat på ett stickprov.  
Syntax  
VARIANS( tal 1; tal 2; ...tal 30)  
tal 1, tal 2...tal 30 är numeriska argument som utgör ett stickprov från en population.  
Du kan även ange referenser.  
Exempel  
=VARIANS( A1:A50)  
MEDELAVV, MEDEL, TYPVÄRDE, STDAV  
VARIANSA  
Beräknar en uppskattning av variansen baserat på ett stickprov.  
Text värderas till 0.  
Syntax  
VARIANSA( värde 1; värde 2; ...värde 30)  
värde 1, värde 2...värde 30 är argument som utgör ett stickprov ur en population.  
Du kan även ange referenser.  
Text värderas därvid till 0.  
Exempel  
=VARIANSA( A1:A50)  
VARIANS, STDAV och STDAVA  
VARIANSP  
Beräknar variansen baserat på populationen.  
Syntax  
VARIANSP( tal 1; tal 2; ...tal 30)  
tal 1, tal 2...tal 30 är numeriska argument som utgör en population.  
Exempel  
=VARIANSP( A1:A50)  
MEDELAVV, MEDEL, TYPVÄRDE, STDAVP  
VARIANSPA  
Beräknar variansen baserad på populationen.  
Text värderas till 0.  
Syntax  
VARIANSPA( värde 1; värde 2; ...värde 30)  
värde 1, värde 2...värde 30 är argument som utgör en population.  
Exempel  
=VARIANSPA( A1:A50)  
STDAVP och STDAVPA  
PERMUT  
Beräknar antalet möjligheter att dra k element ur en mängd av n element utan upprepning.  
Syntax  
PERMUT( antal_1; antal_2)  
antal_1 är det totala antalet element.  
antal_2 är antalet dragna element.  
Exempel  
=PERMUT( 6; 3) returnerar 120.  
Det finns 120 olika möjligheter att bland 6 spelkort dra en följd av 3 kort.  
BINOMFÖRD, FAKULTET, HYPGEOMFÖRD, KOMBIN, KRITBINOM, NEGBINOMFÖRD  
PERMUT2  
Beräknar antalet möjligheter att dra k element ur en mängd av n element när det dragna elementet läggs tillbaka efter varje dragning.  
Syntax  
PERMUT2( antal_1; antal_2)  
antal_1 är det totala antalet element.  
antal_2 är antalet dragna element.  
Exempel  
Hur många olika kombinationer av 2 element kan göras i en uppsättning av 11 element?  
PERMUT2( 11;2) returnerar 121.  
PERMUT2( 6; 3) returnerar 216.  
Det finns 216 olika möjligheter att bland 6 spelkort dra en följd av 3 kort om Du lägger tillbaka varje draget kort igen innan Du drar nästa.  
BINOMFÖRD, FAKULTET, HYPGEOMFÖRD, KOMBIN2, KRITBINOM, NEGBINOMFÖRD  
SANNOLIKHET  
Beräknar sannolikheten för ett slutet intervall begränsat av två värden.  
Om Du inte anger någon övre gräns, beräknas sannolikhetsfunktionen under antagandet av att de värden som hör till data är lika med det undre gränsvärdet.  
Syntax  
SANNOLIKHET( data; sannolikheter; start; slut)  
data är matrisen med data i stickprovet.  
sannolikheter är matrisen för de tillhörande sannolikheterna.  
start är starten på värdeintervallet vars sannolikheter ska summeras.  
slut (valfritt) är slutet på värdeintervallet vars sannolikheter ska summeras.  
Om denna parameter saknas, beräknas sannolikheten för värdet start.  
Exempel  
=SANNOLIKHET( A1:A50; B1:B50; 50; 60) beräknar sannolikheten för att ett värde i området A1:A50 ligger innanför gränserna 50 och 60.  
För varje värde i området A1:A50 finns en tillhörande sannolikhet i området B1:B50.  
BINOMFÖRD, KRITBINOM  
WEIBULL  
Beräknar sannolikheten för en Weibull-fördelad slumpvariabel.  
Syntax  
WEIBULL( tal; alfa; beta; K)  
tal är värdet för vilket Weibull-fördelningen ska beräknas.  
alfa är Weibull-fördelningens alfa-parameter.  
beta är Weibull-fördelningens beta-parameter.  
K är funktionstypen.  
Om K= 0 beräknas täthetsfunktionen; om K=1 beräknas fördelningen.  
Exempel  
=WEIBULL( 2; 1; 1; 1) returnerar 0,86.  
EXPONFÖRD  
Operatorer i %PRODUCTNAME Calc  
I %PRODUCTNAME Calc kan du använda följande operatorer.  
Aritmetiska operatorer  
Dessa operatorer ger numeriska resultat.  
Operator  
Namn  
Exempel  
+ (plus)  
Addition  
1+1  
- (minus)  
Subtraktion  
2-1  
- (minus)  
Negation  
-5  
* (asterisk)  
Multiplikation  
2*2  
/ (snedstreck)  
Division  
9 / 3  
% (procent)  
Procent  
15%  
^ (inskjutningstecken)  
Exponent  
3^2  
Relationsoperatorer  
Dessa operatorer ger det logiska värdet SANT eller FALSKT.  
Operator  
Namn  
Exempel  
= (likhetstecken)  
Lika med  
A1=B1  
> (större än)  
Större än  
A1>B1  
< (mindre än)  
Mindre än  
A1<B1  
>= (större än eller lika med)  
Större än eller lika med  
A1>=B1  
<= (mindre än eller lika med)  
Mindre än eller lika med  
A1<=B1  
<> (inte lika med)  
Inte lika med  
A1<>B1  
Textoperator  
Operatorn länkar enskilda texter till en hel text.  
Operator  
Namn  
Exempel  
& (och)  
Textoperator Och  
"Sun" & "day "returnerar "Sunday"  
Referensoperatorer  
Dessa operatorer länkar cellområden.  
Operator  
Namn  
Exempel  
: (kolon)  
Område  
A1:C108  
! (utropstecken)  
Snitt  
SUMMA( A1:B6!B5:C12)  
Här ligger cellerna B5 och B6 i snittet och deras summa beräknas.  
Namn  
Med detta kommando kan du definiera namn för de olika områdena i tabellerna.  
Att tilldela områdesnamn gör det lättare att navigera genom tabelldokument och att hitta det man söker.  
Definiera...  
Klistra in...  
Överta...  
Etiketter...  
Definiera namn  
Här kan du ange ett namn på ett cellområde eller på formler och delar av formler.  
Du kan definiera områden med musen eller genom att mata in referensen i inmatningsfälten.  
I kombinationsfältet Tabellområde till vänster på formellisten finns en lista över områdenas namn.  
Motsvarande område i tabellen markeras då.  
Namn som du har definierat för formler eller delar av formler finns inte med här.  
Namn  
Gå till textfältet och skriv namnet på det område eller den formel respektive formeldel som Du vill definiera i det aktuella tabelldokumentet.  
Listrutan ger en överblick över alla de namn som redan är definierade.  
Om Du klickar på ett namn på listan, markeras tillhörande områdeshänvisning i dokumentet med en blå ram.  
Om flera cellområden hör till samma områdesnamn, visas de samtidigt i avvikande färg.  
Hänvisar till  
Här anger Du en områdeshänvisning för det valda områdesnamnet, eller också för Du in en formel, t ex =A1+1 eller $A1*20, som Du vill kunna hänvisa till med det valda namnet.  
Om Du vill mata in en ny områdeshänvisning, kan Du placera insättningspunkten i det här fältet och direkt föra in hänvisningen genom att markera tabellområdet i fråga på det aktuella bladet eller på ett annat blad.  
Fler  
Välj den här kommandoknappen när Du vill utvidga namngivningen med tillägget Typ av område.  
Typ av område  
Här kan Du ange områdestyp för den valda områdesdefinitionen.  
Utskriftsområde  
Om Du vill definiera områdesdefinitionen som ett utskriftsområde, klickar Du här.  
Filter  
Här kan Du definiera den valda områdesdefinitionen som filter.  
Upprepningskolumn  
Här kan Du definiera den valda områdesdefinitionen som upprepningskolumn.  
Upprepningsrad  
Här kan Du definiera den valda områdesdefinitionen som upprepningsrad.  
Fler  
Med den här kommandoknappen stänger du tilläggsområdet.  
Lägg till / Ändra  
Med kommandoknappen Lägg till lägger du till ett nytt namn i namnlistan, och med Ändra kan du ändra ett redan angivet namn som du väljer på namnlistan.  
Infoga namn  
Här väljer Du ett tidigare definierat cellområde som ska infogas där markören står i dokumentet.  
Detta görs genom att Du markerar områdesnamnet.  
Du kan inte infoga ett namn om Du inte tidigare har gett området namnet.  
Infoga namn  
Här visas en förteckning över de döpta områdena i tabellen.  
Om Du dubbelklickar på en post, infogas motsvarande område i tabellen där markören står.  
Lista  
Här infogar Du en lista över cellreferenserna till alla de döpta områden där markören står i tabellen.  
Skapa namn  
I den här dialogrutan bestämmer du att namn för markerade cellområden ska skapas automatiskt.  
Markera först alla de celler som ska få ett namn som område.  
Därefter öppnar du den här dialogrutan.  
Skapa namn från  
I detta område kan Du bestämma ur vilken del av tabellen namnet ska skapas.  
Sidhuvud  
Om Du vill skapa områdesnamn ur posterna i det markerade tabellområdets första rad klickar Du här.  
Varje kolumn får ett separat namn och en cellreferens.  
Vänstra kolumnen  
Här kan Du skapa områdesnamn ur posterna i den första kolumnen i det markerade tabellområdet.  
Varje rad får ett separat namn och en cellreferens.  
Sidfot  
Om Du vill skapa områdesnamn ur posterna på det markerade tabellområdets sista rad klickar Du här.  
Varje kolumn får ett separat namn och en cellreferens.  
Högra kolumnen  
Här kan Du skapa områdesnamn ur posterna i den sista kolumnen i det markerade tabellområdet.  
Varje rad får ett separat namn och en cellreferens.  
Definiera etikettområde  
I den här dialogrutan definierar du ett etikettområde.  
Det enskilda innehållet i cellerna i ett etikettområde kan du infoga som namn i formler - %PRODUCTNAME känner sedan igen dessa namn på samma sätt som t.ex. de fördefinierade namnen på veckodagar och månader.  
Det betyder att namnet kompletteras automatiskt vid inmatning i en formel.  
Dessutom har etikettområdena högre prioritet än automatiskt skapade områden om ett namn skulle förekomma flera gånger.  
Du kan definiera flera etikettområden som innehåller samma etiketter på olika tabeller.  
I sådana fall kontrollerar %PRODUCTNAME först den aktuella tabellens områden och, om sökningen inte ger något resultat, kontrolleras därefter övriga tabellers områden.  
Område  
Här visas varje etikettområdes cellområde.  
Om du vill radera ett etikettområde igen, markerar du det och klickar sedan på Radera.  
innehåller kolumnhuvuden  
Välj det här alternativet om det aktuella etikettområdet ska innehålla kolumnhuvuden.  
innehåller radhuvuden  
Välj det här alternativet om det aktuella etikettområdet ska innehålla radhuvuden.  
för dataområde  
I det här textfältet visas det definierade tabellområdet.  
Du kan ändra området när dialogrutan har öppnats genom att klicka i tabellen och välja ut ett annat område genom att markera det med musen.  
Lägg till  
Här läggs det aktuella etikettområdet till i listan.  
Funktioner  
Med det här kommandot öppnar du funktionsfönstret, där du har tillgång till samtliga funktioner som du kan infoga i dokumentet.  
Funktionsfönstret är ett förankringsbart fönster vars storlek du kan ändra.  
Med dess hjälp kan du snabbt mata in funktioner i tabelldokumentet.  
När du dubbelklickar på en post i funktionslistan infogas motsvarande funktion direkt med alla parametrar.  
Kategorilista  
Funktionslista  
I den här listrutan listas de funktioner som tillhör den valda kategorin.  
Välj ut den önskade funktionen med musen.  
När Du klickar på någon funktion visas en kort funktionsbeskrivning i funktionsfönstrets nedre del.  
Om Du vill infoga den markerade funktionen i dokumentet dubbelklickar Du på den eller på ikonen Infoga funktion i beräkningsark.  
Infoga funktion i beräkningsark  
Om du klickar på den här ikonen infogas den markerade funktionen i dokumentet.  
Här öppnar du en dialogruta där du kan välja ut en fil.  
Externa data  
Här infogar du externa data (webbsidessökningar) i en tabell.  
URL för extern datakälla  
Ange från vilken URL eller fil som de externa data laddas.  
Tillgängliga tabeller / områden  
Här väljer du ett område eller en tabell.  
Uppdatering var  
Här definierar du hur ofta externa data ska laddas om och visas.  
Cellattribut  
Med det här kommandot kan du välja olika formatalternativ och tilldela de markerade cellerna.  
Tal  
Teckensnitt  
Cellskydd  
Här kan du förse markerade celler med olika skyddsalternativ.  
Skydd  
I det här området kan du välja mellan skyddsalternativen Skyddad, Dölj formel och Dölj allt.  
Skyddad  
Om du vill skydda de markerade cellerna mot förändringar klickar du här.  
Detta cellskydd fungerar bara om du även skyddar tabellen (Verktyg - Skydda dokument - Tabell).  
Dölj formel  
Här kan du definiera att formlerna i de markerade cellerna ska döljas.  
Dölj allt  
Om du väljer det här alternativet döljs formler och innehåll i de markerade cellerna.  
Utskrift  
Här kan du göra standardinställningar för hur din tabell ska skrivas ut.  
Dölj vid utskrift  
Om du aktiverar det här fältet skrivs de markerade cellerna inte ut.  
Rad  
Med här undermenyerna kan du ställa in radhöjd och dölja eller visa markerade rader.  
Höjd...  
Optimal höjd...  
Optimal radhöjd  
Här väljer du den optimala radhöjden för de markerade raderna.  
Du kan använda olika måttenheter i %PRODUCTNAME Calc.  
Extra  
Med det här rotationsfältet definierar du ett ytterligare avstånd mellan det största tecknet på en rad och cellavgränsningarna.  
Standardvärde  
Återställer standardvärdet för den optimala radhöjden.  
Det ytterligare avståndet för den optimala radhöjden sätts till 0,0 cm.  
Dölj  
Med det här kommandot döljer du markerade rader, kolumner eller tabeller.  
Kolumn - Dölj.  
Du kan dölja en enskild tabell genom att klicka på den aktuella tabellfliken och sedan välja kommandot Format - Tabell - Dölj.  
Dolda tabeller skrivs inte ut om de inte ingår i ett utskriftsområde.  
Om det finns dolda rader eller kolumner visas de som avbrott i rad - / kolumnhuvudena.  
Om du vill visa dolda rader, kolumner eller tabeller igen väljer du Format - Rad / Kolumn - Visa eller Format - Tabell - Visa.  
Visa  
Med det här kommandot kan du visa dolda rader eller kolumner igen.  
Om Du vill visa rader eller kolumner, markera ett område med rader eller kolumner, som omger de dolda elementen, och välj kommandot Format - Rad - Visa eller Format - Kolumn - Visa.  
Kolumn  
Här hittar du undermenykommandona med vilka du ställer in kolumnbredd och visar och döljer kolumner.  
Bredd...  
Optimal bredd...  
Optimal kolumnbredd  
Här väljer du den optimala kolumnbredden för de markerade kolumnerna.  
Du kan använda olika måttenheter i %PRODUCTNAME Calc.  
Extra  
Med hjälp av det här rotationsfältet definierar du ett ytterligare avstånd mellan den längsta posten i en kolumn och de vertikala kolumnkanterna.  
Standardvärde  
Med det här alternativet ställer du in den optimala kolumnbredd med vilken hela kolumnens innehåll visas, utan att texten "rinner ut" ur kolumnen.  
Det extra avståndet för den optimala kolumnbredden sätts till 0,2 cm.  
Tabell  
Med det här kommandot öppnar du en undermeny, där du kan byta namn på den aktuella tabellen och dölja den.  
Om du redan har dolt en tabell öppnas en dialogruta, där du kan välja en tabell som ska visas igen.  
Byt namn...  
Visa...  
Byt namn  
En dialogruta öppnas där du kan ge den aktuella tabellen / kalkylarket ett annat namn.  
Namn  
I det här textfältet anger du tabellens / kalkylarkets namn.  
Du kan också öppna den här dialogrutan via den snabbmeny som visas om du trycker på musknappen tillsammans med Ctrl-tangenten högra musknappen i tabellfliksområdet i fönstrets nederkant.  
Du kan även klicka på tabellfliken och samtidigt hålla ner Kommando Alt -tangenten.  
Nu kan du ändra namnet direkt.  
Visa tabell  
Med det här kommandot kan du åter visa tabeller som har dolts med kommandot Dölj.  
Bara en enda tabell får vara markerad, annars går det inte att välja kommandot.  
Den aktuella tabellen är alltid markerad.  
Du avmarkerar en annan tabell genom att klicka på tabellnamnet i den undre fönsterkanten med nedtryckt Kommando Ctrl -tangent.  
Dolda tabeller  
Här visas namnen på de dolda tabellerna.  
Om du vill visa en viss tabell igen, klickar du på en post i listan och bekräftar valet med OK.  
Sammanfoga celler  
Här ser du en undermeny där du kan sammanfoga celler till en gemensam cell och upphäva denna sammanfogning.  
Definiera  
Med det här kommandot sammanfogas det markerade cellområdet, d.v.s. det behandlas som en cell.  
Den sammanfogade cellen får samma celladress som den första cellen i det ursprungliga cellområdet.  
Sammanfogade celler kan inte sammanfogas en gång till med andra celler.  
Området måste vara en rektangel; multipla markeringar stöds inte.  
Om det finns något innehåll i cellerna som ska sammanfogas, så visas en säkerhetskontroll.  
Upphäv  
Med det här kommandot upphäver du sammanfogningen av ett cellområde.  
Välj ut den sammanfogade cellen och välj det här kommandot.  
Sidformatmall  
Med det här kommandot öppnar du en dialogruta där du kan styra utseendet för hela sidor.  
Tabell  
Du anger även ordningsföljden för de utskrivna sidorna, det första sidnumret och skalningen här.  
Skriv ut  
I det här området bestämmer du vilka tabellelement som ska skrivas ut.  
Rad - och kolumnhuvuden  
Markera den här rutan om du vill skriva ut kolumnhuvudena A, B,... och radhuvudena 1, 2,... i marginalerna på de utskrivna sidorna.  
Tabellgitter  
Markera här om begränsningarna av de enskilda cellerna i ett gitternät ska skrivas ut.  
Välj Verktyg - Alternativ - Tabelldokument - Vy och markera Gitterlinjer om du vill göra inställningen för vyn på bildskärmen.  
Anteckningar  
Markera den här rutan om du vill skriva ut anteckningarna i tabellen.  
De hamnar på en egen sida, och framför varje anteckning anges adressen till motsvarande cell.  
Objekt / grafik  
Om du har markerat den här rutan, skrivs även infogade objekt (om de kan skrivas ut) och grafikobjekt ut.  
Diagram  
Markera det här alternativet om du vill skriva ut integrerade diagram.  
Ritobjekt  
Om du markerar den här rutan, skrivs de objekt som du själv har ritat ut.  
Formler  
Markera det här fältet när du vill skriva ut formlerna i stället för de uträknade resultaten.  
Nollvärden  
Markera den här rutan om talet 0 ska skrivas ut.  
I annat fall skrivs celler med värdet Noll inte ut.  
Sidordning  
Här definierar du ordningsföljden som ska gälla när flersidiga tabeller ska delas upp på de utskrivna sidorna.  
Uppifrån och ned  
Markera det här alternativet om du vill att de vänstra kolumnerna fram till tabellens nederkant ska skrivas ut först.  
Från vänster till höger  
Markera det här alternativet om du vill att de övre raderna fram till tabellens högerkant ska skrivas ut först.  
Första sidnummer  
Markera det här fältet om du vill ange ett annat första sidnummer än 1.  
Den första sidan får det sidnummer som du har ställt in i rotationsfältet.  
Skalning  
I det här området definierar du en skala för utskriften av tabelldokument på papper.  
Förminska / förstora utskrift  
Om du markerar det här alternativet, kan du i rotationsfältet till höger välja en förstorings - eller förminskningsfaktor som alla utskrivna sidor ska skalas med.  
Mata in skalningsfaktorn här.  
Anpassa utskrift till antal sidor  
Om du markerar det här alternativet kan du i rotationsfältet till höger ange ett maximalt antal utskriftssidor som hela dokumentet ska skrivas ut på.  
Det skalas då så att det får rum på de sidorna.  
Mata in det maximala antalet sidor som ska skrivas ut här.  
Utskriftsområden  
Här kan du definiera ett utskriftsområde för varje tabell för sig.  
Om du har definierat ett utskriftsområde skrivs bara det definierade utskriftsområdet ut när tabellen skrivs ut.  
Du kan dessutom ange att en viss rad eller kolumn ska skrivas ut på varje följande sida.  
Redigera...  
Definiera  
Med det här kommandot kan du definiera en aktiverad cell eller ett markerat, sammanhängande cellområde som utskriftsområde.  
Upphäv  
Med det här kommandot kan du upphäva ett utskriftsområde som har definierats för den aktuella tabellen.  
Redigera utskriftsområden  
Med det här kommandot öppnar Du en dialogruta, där Du kan ange inställningar för utskriftsområdet.  
Du kan även definiera upprepningsrader eller upprepningskolumner, som ska skrivas ut på varje sida.  
Utskriftsområde  
Här kan Du ange inställningar för ett definierat utskriftsområde.  
I kombinationsrutan väljer Du ett definierat utskriftsområde.  
Välj -ingen - om Du vill upphäva ett definierat utskriftsområde i den aktuella tabellen.  
Välj -markering - om Du vill definiera det markerade området i tabellen som utskriftsområde.  
Med -användardefinierad - kan Du ange ett utskriftsområde som Du tidigare har definierat med kommandot Format - Utskriftsområden - Definiera.  
Om Du t ex har namngett ett område med Infoga - Namn - Definiera så visas namnet i listrutan, i vilken Du kan välja det.  
I textrutan till höger kan Du ange ett utskriftsområde med cellreferenser eller som områdesnamn.  
När markören i står i textrutan Utskriftsområde kan Du även markera ett utskriftsområde i tabellen med musen.  
Upprepningsrad  
Här kan Du välja en eller flera rader, som ska upprepas på varje sida vid utskrift.  
I textrutan till höger anger Du en radreferens enligt mönstret "1" eller "$1 "eller "$2:$3".  
I kombinationsrutan visas då -användardefinierad -.  
Om Du väljer -inga - upphävs den definierade upprepningsraden.  
Du kan även definiera upprepningsrad( er) genom att dra med musen i tabellen när markören står i textfältet Upprepningsrad.  
Upprepningskolumn  
Här kan Du välja en eller flera kolumner, som ska upprepas på varje sida vid utskrift.  
I textrutan till höger anger Du en kolumnreferens enligt mönstret "A", "AB", "$A" eller "$C:$E ".  
I kombinationsrutan visas då -användardefinierad -.  
Om Du väljer -inga - upphävs den definierade upprepningskolumnen.  
Du kan även definiera upprepningskolumn( er) genom att dra med musen i tabellen när markören står i textfältet Upprepningskolumn.  
Lägg till  
Med det här kommandot lägger du till den aktuella markeringen till de utskriftsområden som har definierats för tabellen.  
Mallkatalog  
Med det här alternativet öppnar du mallkatalogen där du kan skapa, redigera och administrera formatmallar och dokumentmallar.  
Förutom administrationen av mallar har Stylist samma funktioner.  
Malltyp  
I det här kombinationsfältet anger du om cell - eller sidformatmallar ska visas i mallförteckningen.  
Mallista  
Här visas en lista med mallarna i det valda mallområdet.  
På snabbmenyn kan du välja kommandon för att skapa en ny mall, radera en egen mall eller ändra den markerade mallen.  
Mallområde  
De färdiga mallarna är uppdelade i flera formatmallsområden så att förteckningen ska bli överskådlig.  
Alla mallar  
Visar alla mallar för den aktuella malltypen.  
Använda mallar  
De är också tillgängliga på objektlisten.  
Användardefinierade formatmallar  
Visar de formatmallar av den aktuella typen som har definierats av någon användare.  
Hierarkiskt  
Visar formatmallarna av den aktuella typen i hierarkisk uppställning.  
Den här uppställningen liknar mallstrukturen på hårddisken.  
Om Du vill se mallarna på nivån under, klickar Du på plustecknet intill mallnamnet.  
Nytt...  
Välj det här kommandot om du vill skapa en ny mall.  
Beroende på malltyp öppnas dialogrutan Cellformatmall eller Sidformatmall.  
Ändra...  
Välj det här kommandot om Du vill ändra den markerade mallen.  
Beroende på malltyp öppnas dialogrutan Cellformatmall eller Sidformatmall.  
Radera...  
Välj det här kommandot om du vill radera den markerade mallen.  
Du kan bara radera användardefinierade formatmallar.  
Innan raderingen utförs ombeds du bekräfta den.  
Administrera...  
När du klickar på den här kommandoknappen öppnas dialogrutan för administration av dokumentmallar.  
Stylist  
Med det här kommandot visar och döljer du Stylist.  
Med Stylist tilldelar du objekt och textområden formatmallar.  
Du kan uppdatera objekt och textområden, ändra existerande mallar och skapa nya mallar.  
Du kan låta det förankringsbara fönstret vara öppet medan du redigerar dokumentet.  
Cellformatmallar  
Här väljer du listan över cellformatmallarna för indirekt formatering av celler.  
Cellformatmallar  
Sidformatmallar  
Här väljer du listan över sidformatmallar för indirekt formatering av sidlayouten.  
Sidformatmallar  
Tilldelningsläge  
Sätter på och stänger av tilldelningsläget.  
I det här läget tilldelar du den mall som har markerats i Stylist.  
Tilldelningsläge  
Så här tilldelar du en ny formatmall i tilldelningsläget:  
Markera en mall i Stylist.  
Klicka på ikonen Tilldelningsläge.  
Flytta muspekaren till det objekt eller det område som du vill tilldela den aktuella formatmallen.  
Tryck ned den vänstra musknappen om Du vill formatera en cell, eller dra med nedtryckt musknapp över flera celler för att formatera dem alla.  
Upprepa vid behov den här proceduren för ytterligare celler och områden.  
Klicka på nytt på ikonen Tilldelningsläge om du vill avsluta det här läget.  
Ny formatmall av markering  
Här skapar du en ny mall som innehåller formateringen av det markerade objektet.  
Du döper den nya formatmallen i dialogrutan Skapa formatmall som visas automatiskt.  
Skapa ny formatmall av markering  
Uppdatera formatmall  
Här övertar den mall, som har markerats i Stylist, den aktuella formateringen av det markerade objektet.  
Uppdatera formatmallar  
Snabbmenyn - Nytt... / Ändra... / Radera...  
Här har Du tillgång till samma funktioner som i dialogrutan Format - Mallkatalog.  
Mallkategori  
I det här kombinationsfältet väljer du en mallkategori.  
AutoFormat  
Med det här kommandot kan du tilldela ett markerat tabellområde ett AutoFormat och definiera egna AutoFormat.  
Fr.o.m. version %PRODUCTNAME 5.0 kan Du även överta roterade texter till AutoFormat och använda dem som AutoFormat.  
Detta innebär att det filformat som används för att spara AutoFormat i %PRODUCTNAME Writer och %PRODUCTNAME Calc är inkompatibelt med tidigare versioner. %PRODUCTNAME 5.0, 5.1 och %PRODUCTVERSION kan fortfarande läsa det gamla formatet, men äldre versioner av %PRODUCTNAME kan inte läsa det nya AutoFormatet.  
Cellformat  
Du kan välja ut något av dessa AutoFormat och tilldela det markerade tabellområdet AutoFormatet.  
Lägg till...  
Klicka på Lägg till.  
Ange ett namn och klicka på OK.  
Fler >>  
Med denna kommandoknapp öppnar Du området Formatering, där Du kan utesluta enstaka formateringsalternativ i AutoFormat.  
Formatering  
I det här området kan Du utöka dialogrutan AutoFormat med alternativen Talformat, Inramning, Teckensnitt, Mönster, Justering och Anpassa bredd och höjd.  
Talformat  
Avmarkera kryssrutan om talformatet inte ska ändras.  
Inramning  
Avmarkera om inramningen inte ska ändras.  
Teckensnitt  
Avmarkera om teckensnittet inte ska ändras.  
Mönster  
Avmarkera om mönstret (färger, etc) inte ska ändras.  
Justering  
Avmarkera om justeringen inte ska ändras.  
Anpassa bredd och höjd  
Avmarkera om bredden och höjden inte ska ändras.  
Byt namn  
Klicka på den här kommandoknappen om Du vill ändra beteckningen på det valda AutoFormatet.  
Kommandoknappen är bara synlig om Du har valt Fler >>.  
Dialogen Byt namn på AutoFormat öppnas.  
Mata in det nya namnet på AutoFormatet här.  
Fler <<  
Med den här kommandoknappen döljer Du tilläggsalternativen i området Formatering.  
Villkorlig formatering  
I dialogrutan Villkorlig formatering kan du definiera formatmallar beroende på villkor.  
Om en cell redan tilldelats en formatmall ändras denna aldrig.  
För den formatmall som du anger här görs då en extra utvärdering.  
Du kan ange upp till tre villkor som antingen söker på innehållet i cellvärden eller i formler.  
Sökning på villkoren sker i tur och ordning från villkor 1 till villkor 3.  
I annat fall sker sökning på villkor 2 och om det uppfylls används formatmallen för detta.  
Om villkor 2 inte uppfylls sker även sökning på villkor 3.  
Bland exemplen för %PRODUCTNAME finns dokumentet {installpath} / share / samples / swedish / spreadsheets / biorytm.sdc, där villkorlig formatering använts i tabellen "Detaljer ".  
Villkor 1 / 2/3  
Markera den här rutan om du vill definiera ett villkor.  
För varje villkor markerar du respektive ruta och sedan skriver du in villkoren.  
Du stänger dialogrutan med OK.  
Cellvärde / Formel  
I det här kombinationsfältet väljer du om den villkorliga formateringen ska vara beroende av ett cellvärde eller en formel.  
Om du väljer en formel som referens döljs kombinationsfältet Cellvärdesvillkor direkt till höger om fältet Cellvärde / Formel.  
Om den aktuella cellen innehåller ett värde som inte är lika med noll så uppfylls villkoret.  
Cellvärdesvillkor  
Om detta villkor uppfylls formateras de markerade cellerna enligt den definierade formatmallen.  
I kombinationsfältet Cellvärdesvillkor, som bara visas om du kontrollerar ett cellvärde, väljer du ett villkor för att de markerade cellerna ska formateras enligt den definierade formatmallen.  
Om du har valt ett villkor som kräver två parametrar (t.ex. "mellan "eller "inte mellan"), delas parameterfältet in i två parameterfält med varsin Förminska - / Förstora-ikon.  
Cellformatmall  
Här väljer du mallen som ska användas när villkoret uppfylls.  
Parameterfält  
Här anger du en referens, ett värde eller en formel.  
Du anger en referens, ett värde eller en formel i parameterfältet (eller i de två parameterfälten, om du har valt ett villkor som kräver två parametrar).  
Du kan även använda formler med relativa referenser.  
På det här sättet kompletteras villkoret.  
Det kan t.ex. se ut så här:  
Cellvärdet är lika med 0:  
Cellformatmall Nollvärde (exemplet förutsätter att du har definierat en cellformatmall med namnet Nollvärde, som ska framhäva nollvärden).  
Cellvärdet är mellan $B$20 och $B$21:  
Cellformatmall Resultat (exemplet förutsätter att aktuella gränsvärden finns angivna i cellerna B20 och B21 samt att cellformatmallen Resultat finns).  
Formeln är SUMMA( $A$1:$A$5 )=10:  
Cellformatmall Resultat (de markerade cellerna formateras enligt formatmallen Resultat om summan av innehållet i cell A1 t o m A5 är lika med 10).  
Cellformatmall  
Här kan du skapa en cellformatmall.  
Tal  
Avstavning  
Det här menykommandot öppnar dialogrutan där du kan ställa in avstavningen i %PRODUCTNAME Calc.  
Du kan bara använda den automatiska avstavningen i %PRODUCTNAME Calc om Radbrytning är aktiverad.  
Avstavning för markerade celler  
Markera cellerna där du vill ändra avstavningen.  
Välj kommandot Verktyg - Avstavning.  
Dialogrutan Cellattribut öppnas med fliken Justering.  
Markera rutan Avstavning aktiv.  
Avstavning för ritobjekt  
Markera ett ritobjekt.  
Välj kommandot Verktyg - Avstavning.  
Varje gång du väljer kommandot sätter du på eller stänger av avstavningen för ritobjektet.  
En bock visar aktuell status.  
Detektiv  
Med det här kommandot öppnar du tabelldokument-detektiven.  
Med hjälp av detektiven kan du synliggöra sambanden mellan den aktuella formelcellen och andra celler i tabellen.  
Om du har definierat ett spår i tabellen kan du föra markören till spåret.  
Den förvandlas då till ett förstoringsglas med hänvisningspilar.  
Om du dubbelklickar med den här markören på det synliga spåret så markeras cellen i bortre änden av spåret.  
Spår till överordnade  
Denna funktion visar spåret mellan den aktuella formelcellen och cellerna som används i formeln.  
Spår i tabellen visas med markeringspilar Samtidigt framhävs området med alla celler som används i formeln i den aktuella cellen med en blå ram.  
Funktionen arbetar nivå för nivå.  
Om t.ex. spåret från en formel till dess överordnade celler redan visas, skapas spåren till deras överordnade celler i sin tur om funktionen används igen.  
Ta bort spår till överordnade  
Den här funktionen raderar en nivå med markeringspilar som infogats med Spår till underordnade.  
Spår till underordnade  
Den här funktionen skapar markeringspilar från den aktuella cellen till formelcellerna som använder värdet i den aktuella cellen.  
Samtidigt framhävs området med alla celler som används tillsammans med den aktuella cellen i en formel med en blå ram.  
Funktionen arbetar nivå för nivå.  
När t.ex. spåret från en cell till dess underordnade cell (t.ex. formeln som använder den här cellen som referens) redan visas, skapas i sin tur spåren till deras underordnade celler nästa gång du använder funktionen.  
Ta bort spår till underordnade  
Den här funktionen raderar en nivå med markeringspilarna som har infogats med Spår till underordnade.  
Ta bort alla spår  
Med detta kommando tar du bort alla markeringspilar (spår) som infogats med Detektiv i tabellen.  
Spår till fel  
Den här funktionen visar de överordnade cellerna till en markerad cell som innehåller en felkod.  
Fyllningsläge  
Med den här funktionen aktiverar du detektivens fyllningsläge.  
Muspekaren förvandlas till en fyllningsläge-ikon, och du kan titta på spåren till överordnade celler från valfria celler som du klickar på.  
Du avslutar det här läget genom att trycka på Esc-tangenten eller välja kommandot Avsluta fyllningsläge på snabbmenyn.  
Funktionen Fyllningsläge är identisk med kommandot Spår till överordnade när den aktiveras första gången.  
På snabbmenyn kan du välja fler alternativ för fyllningsläget och avsluta fyllningsläget.  
Ringa in ogiltiga data  
Med den här funktionen ringar du in cellerna i tabellen vars innehåll inte motsvarar giltighetsreglerna.  
Med giltighetsregler kan du vid behov begränsa inmatningen av tal, datum, tider och texter till vissa värden.  
Med det är ändå möjligt att mata in ogiltiga värden (så länge du inte har valt åtgärden "Stopp") eller att kopiera ogiltiga värden till cellerna.  
Dessutom ändras inte värden som finns i celler om du först i efterhand tilldelar en giltighetsregel.  
Uppdatera spår  
Med det här kommandot uppdaterar du de visade spåren.  
Då tas formler som eventuellt har ändrats under tiden med vid visning av spåren.  
Detektiv-pilar i dokumentet uppdateras om följande villkor uppfylls:  
Om du har valt Verktyg - Detektiv - Uppdatera spår.  
Om du har aktiverat alternativet Verktyg - Detektiv - Uppdatera automatiskt för varje ändring av formler i dokumentet.  
Uppdatera automatiskt  
Med denna omkopplare anger du att Detektiv-pilarna ska uppdateras automatiskt så snart en formel ändras.  
Målvärdessökning  
Med det här kommandot öppnar du en dialogruta, där du kan lösa ekvationer med en variabel.  
När sökningen är färdig visas resultatet i en dialogruta.  
Du kan använda resultatet och målvärdet i din beräkning.  
Förinställningar  
I det här området definierar du variablerna.  
Formelcell  
Formelcellen innehåller adressen till den cell där formeln har lagts in.  
Den aktuella celladressen visas redan där.  
Om du klickar på en annan cell i tabellen infogas en referens till den i textrutan.  
Målvärde  
Här anger du målvärdet, d.v.s. svaret på frågeställningen.  
Variabel cell  
I det här fältet läggs celladressen in.  
Den innehåller ett föränderligt värde.  
Skapa scenario  
Här kan du definiera ett scenario för det markerade tabellområdet.  
Namn på scenariot  
Här kan du ange eller ändra namnet för scenariot (på snabbmenyn Egenskaper... i Navigator).  
Du väljer nämligen vy (och senare redigering) för scenarier utifrån det namn som visas på tabellflikarna i fönstrets undre kant eller i Navigator.  
Kommentar  
Här kan du ange eller ändra ytterligare kommentarer till scenariot (på snabbmenyn Egenskaper... i Navigator).  
Kommentarerna visas i Navigator om du klickar på ikonen Scenarion och väljer ett scenario.  
Inställningar  
I det här området gör du inställningar för hur scenarierna ska visas.  
Visa ram  
Du väljer ramens färg i kombinationsfältet.  
Ramen innehåller en titellist där namnet på det senaste scenariot visas.  
När du klickar på den visas en översikt över alla scenarier i det här området om du har definierat flera scenarier.  
Från den här listan kan du välja vilket scenario du vill.  
Kopiera tillbaka  
Om du klickar på den här rutan kopieras först data till det aktiva scenariot tillbaka när du väljer ett scenario.  
Du kan sedan redigera data för varje scenario direkt i tabellen.  
Om du inte väljer det här alternativet i kombination med Visa ram visas inga scenarier i tabellen.  
Då kan du bara använda Navigator.  
Tryck på kommandoknappen Scenarion i Navigator så att alla scenarier i tabellen visas och kan väljas.  
Kopiera hel tabell  
Markera den här rutan om du vill att hela tabellen ska kopieras till en särskild scenario-tabell.  
Skydda dokument  
Med det här kommandot kan du skydda tabeller och dokument mot ändringar.  
Dessutom kan du skydda det aktuella området med lösenord.  
Tabell...  
Dokument...  
Skydda tabell  
Där kan du med eller utan lösenord skydda tabellen mot ändringar.  
Om du vill skydda cellerna i tabellen mot ytterligare redigering, måste rutan Skyddad vara markerad under fliken Cellskydd i dialogen Cellattribut som du öppnar via menyn Format - Cell... eller snabbmenyn Formatera celler....  
Du kan även definiera oskyddade celler eller cellområden i en för övrigt skyddad miljö genom att kombinera kommandon på menyerna Verktyg - Skydda dokument - Tabell... och Format - Cell... - Cellskydd (eller på snabbmenyn Formatera celler... - Cellskydd).  
Markera först det "fria" området och öppna sedan fliken Cellskydd på menyn Format - Cell... eller på snabbmenyn Formatera celler.  
Avmarkera kryssrutan Skyddad i området Skydd och klicka på OK.  
Aktivera därefter skyddet för tabellen ¨på menyn Verktyg - Skydda dokument - Tabell....  
Från och med nu kan bara det område som Du har definierat ändras.  
Om Du senare vill omvandla ett "fritt" område till ett skyddat, så markerar Du området och markerar kryssrutan Skyddad på menyn Format - Cell... - Cellskydd eller på motsvarande snabbmeny.  
Då är även det område skyddat som tidigare kunde ändras.  
Skyddet för en tabell omfattar även tabellflikarnas snabbmeny vid den nedre bildkanten.  
Du kan inte välja menykommandona Radera... och Flytta / kopiera....  
Du kan inte ändra en skyddad tabell eller ett skyddat tabellområde förrän skyddet upphävs.  
Om Du vill upphäva skyddet använder Du kommandot Verktyg - Skydda dokument - Tabell... igen.  
Om Du inte har tilldelat något lösenord, så upphävs tabellskyddet direkt.  
Om Du dessutom har skyddat tabellen med ett lösenord, så visas nu dialogrutan Upphäv tabellskydd, där Du måste skriva in lösenordet.  
Först då avlägsnas den markeringsbock som visar skyddet.  
När Du har sparat en tabell med skydd kan Du bara spara den på nytt via menyn Arkiv - Spara som..., vilket minskar risken för att Du skriver över filen av misstag.  
Lösenord (valfritt)  
Om Du vill skydda tabellen mot obehöriga och oavsiktliga ändringar, kan Du skriva in ett lösenord här.  
Ett omfattande skydd för ditt arbete får du genom att kombinera de båda möjligheterna på menyn Verktyg - Skydda dokument med ett lösenord.  
Om du vill förhindra att dokumentet överhuvudtaget kan öppnas, markerar du rutan Spara med lösenord första gången du sparar, och klickar först därefter på kommandoknappen Spara.  
Dialogrutan Mata in lösenord öppnas där du kan skriva in en teckensträng och bekräfta med OK.  
Tänk på att om du glömmer lösenordet innebär det att inte ens du själv kan komma åt dokumentet.  
Skydda dokument  
När du öppnar menyn Verktyg - Skydda dokument - Dokument... visas dialogrutan Skydda dokument, där du kan skydda ett dokument mot ändringar med eller utan lösenord.  
Du kan inte ändra strukturen i ett skyddat tabelldokument förrän skyddet upphävts.  
Varken Radera..., Flytta / kopiera... eller något annat alternativ är tillgängligt.  
Om Du vill upphäva skyddet, välj kommandot Verktyg - Skydda dokument - Dokument... igen.  
Om Du inte lagt in något lösenord upphävs skyddet omedelbart.  
Om Du har lagt in ett lösenord öppnas dialogrutan Upphäv dokumentskydd, där Du måste skriva in lösenordet.  
Då tas bocken, som visar att skyddet är aktiverat, bort.  
Ett skyddat dokument kan Du, efter att det sparats, endast spara på nytt via menyn Arkiv - Spara som... vilket hjälper Dig att undvika oavsiktliga ändringar i filen.  
Lösenord (valfritt)  
Om Du vill skydda dokumentets struktur från obehöriga eller mot oavsiktliga ändringar kan Du skriva in ett lösenord här.  
Om Du kombinerar de båda alternativen på menyn Verktyg - Skydda dokument med ett lösenord får Du ett fullgott skydd för Ditt arbete.  
Om Du vill skydda ett dokument så att ingen annan kan öppna det så ska Du markera alternativet Spara med lösenord och sedan klicka på Spara första gången som Du sparar dokumentet.  
Då öppnas dialogrutan Mata in lösenord, där Du skriver in en lämplig teckensekvens och bekräftar med OK.  
Tänk på att om Du glömmer lösenordet så har Du inte ens själv tillgång till dokumentet.  
Automatisk beräkning  
Med det här kommandot beräknas formler automatiskt på nytt och resultatet korrigeras vid behov.  
Den nya beräkningen sker för alla celler när en cell i tabellen har ändrats.  
Även diagram i tabellen uppdateras.  
När du har markerat detta alternativ så är kommandot Beräkna på nytt (F9) inte aktiverat.  
Beräkna på nytt  
Här kan du göra om beräkningen av den aktiva tabellen omedelbart.  
Använd detta kommando om du har stängt av den automatiska beräkningen eller om du vill kontrollera att du verkligen ser den uppdaterade versionen när du arbetar med mycket stora tabeller.  
Efter beräkningen visas dokumentet på nytt i fönstret.  
Även diagrammen i tabellen uppdateras.  
Alla celler beräknas på nytt om du använder tangentkombinationen Skift+Crtl+F9.  
AutoInmatning  
Med det här kommandot aktiverar och inaktiverar du AutoInmatning.  
AutoInmatning kompletterar automatiskt en teckensträng som du matar in med en teckensträng som börjar med samma tecken och som finns i samma kolumn.  
Hela kolumnen inkluderas, upp till en längd på 2000 celler respektive 200 olika strängar.  
När du matar in formler (inmatningen börjar med ett likhetstecken) och strängen överensstämmer entydigt, så visas en lista över de tio senast använda funktionerna i Funktionsautopiloten, alla definierade områdesnamn, alla databasområdesnamn och innehållet i alla etikettområden.  
Du använder tabbtangenten för att bläddra framåt och Skift+Tabb för att bläddra bakåt i listan som visas som tips-hjälp, under förutsättning att det finns flera poster.  
Om du vill använda posten från tips-hjälpen i dokumentet, så trycker du på Retur.  
AutoInmatningen är versalkänslig.  
Om du t.ex. har skrivit "Summa" i en cell kan du alltså inte skriva "summa "i en cell i samma kolumn - i så fall måste du stänga av AutoInmatningen.  
Om flera poster överensstämmer visas en urvalslista.  
Den här listan öppnar Du för den just redigerade kolumnen med tangenterna Ctrl+D eller med snabbmenykommandot Urvalslista....  
Du bläddrar framåt i listan med tabbtangenten, och bakåt med Skift+Tabb.  
Cellinnehåll  
Här öppnar du en undermeny med kommandon för att beräkna tabeller och aktivera AutoInmatning.  
Dela  
När du aktiverar det här menykommandot delas det aktuella fönstret vid det övre vänstra hörnet av den aktuella cellen.  
Du kan även använda musen när Du vill dela arbetsbladets fönster horisontellt eller vertikalt.  
Dra in detta streck i arbetsbladet.  
En tjock svart linje visar var arbetsbladet delas.  
Ett delat fönster får i varje delområde egna bildrullningslister, i motsats till ett fixerat fönsterområde som inte kan rullas.  
Fixera  
Om du aktiverar det här menykommandot delas tabellen i den övre vänstra hörnan av den aktuella cellen och området uppe till vänster fixeras, d.v.s. det går inte att rulla.  
I den här dialogen definierar du ett databasområde i tabellen.  
Namn  
Här kan du definiera ett nytt databasområde eller välja ett befintligt.  
Ange i textfältet namnet på det databasområde som du vill definiera, eller välj namnet på ett befintligt databasområde i listrutan.  
När du har angett namnet markerar du området i tabellen.  
För databasområden är bara enkla rektangulära områden tillåtna.  
Område  
I det här visningsområdet visas vilket område som är kopplat till det valda databasområdet.  
Det område som du markerade när du öppnade dialogrutan visas som förinställning.  
Om du inte har gjort någon markering, markeras det sammanhängande dataområdet där markören står.  
Ändra / Lägg till  
Här införs det för tillfället definierade databasområdet i listan eller också ändras ett befintligt.  
Fler>>  
Om du klickar på den här kommandoknappen utvidgas dialogrutan med området Alternativ.  
Alternativ  
I det här området bestämmer Du alternativ för databasimporten.  
Innehåller kolumnhuvuden  
Välj detta alternativ om det för tillfället definierade databasområdet innehåller kolumnhuvuden.  
Avmarkera det här alternativet om databasområdet inte innehåller några kolumnhuvuden.  
Infoga / radera celler  
Om Du markerar det här alternativet, övertas de rader och kolumner som har infogats i databasen i efterhand i dokumentet.  
För detta behöver Du sedan bara välja kommandot Uppdatera område på menyn Data.  
Alternativet utvärderas även vid filtrering i ett annat område.  
Behåll formatering  
Om Du klickar på den här kryssrutan säkerställer Du att formateringarna bibehålls.  
Om Du t ex har fetformaterat en kolumn och infogar ytterligare en cell ur databasen i kolumnen (menyn Data - Uppdatera område), visas cellens innehåll också fett.  
Spara inte importerade data  
Däremot sparas en hänvisning till databasen.  
Du sparar diskutrymme.  
Källa:  
Här visas information om databasens ursprung och om eventuella operatorer.  
Fler <<  
Klicka här om Du vill förminska den utvidgade dialogrutan.  
Välj område  
Här väljer du ett definierat databasområde.  
Områden  
Här visas alla databasområden som har definierats i det aktuella dokumentet.  
Klicka på en post i listan om du vill välja ett databasområde.  
När du har stängt dialogrutan med OK är databasområdet markerat i tabellen.  
Sortera  
I den här dialogrutan definierar du kriterierna för en sortering.  
Det markerade tabellområdet sorteras alltid efter rader eller kolumner.  
Om du har definierat ett databasområde märker %PRODUCTNAME det automatiskt när markören står i en cell i området.  
Det går inte att sortera om registrering av ändringar är aktiverad.  
Om markören står utanför ett databasområde så skapas ett namnlöst databasområde som används när kommandot väljs.  
Sorteringskriterier  
Här definierar du sorteringskriterierna.  
Du kan välja sorteringsordning, sorteringsriktning och tabellkolumnen eller -raden som ska sorteras.  
Se till att Du även markerar rubrikerna för de rader och kolumner som ska sorteras.  
Sortera efter  
I denna listruta väljer Du det kännetecken som ska ha högsta prioritet vid sorteringen.  
Stigande  
Om detta alternativ är markerat så sorteras stigande, dvs från A till Ö och från 0 till 9.  
Fallande  
Om Du markerar det här alternativet görs en fallande sortering, dvs från Ö till A och från 9 till 0.  
Sedan efter  
I den här listrutan väljer Du det kännetecken som ska ha näst högsta prioritet vid sorteringen.  
Stigande  
Klicka här om sorteringen ska ske stigande, dvs från A till Ö och från 0 till 9.  
Fallande  
Klicka här om sorteringen ska ske fallande, dvs från Ö till A och från 9 till 0.  
Sedan efter  
I den här listrutan väljer Du det kännetecken som ska ha tredje högsta prioritet vid sorteringen.  
Stigande  
Om Du har markerat det här alternativet görs sorteringen stigande, dvs från A till Ö och från 0 till 9.  
Fallande  
Om Du har markerat det här alternativet görs sorteringen fallande, dvs från Ö till A och från 9 till 0.  
Sortera  
Med ikonerna sorterar du de markerade cellerna stigande eller fallande.  
Sifferfält sorteras efter storlek och textfält efter ASCII-ordningsföljden för de tecken som fältet innehåller.  
Ikoner på verktygslisten:  
Alternativ  
Här väljer du alternativen för sorteringen som du har definierat under Sorteringskriterier.  
Versalkänslig  
Om du markerar den här rutan, görs skillnad mellan stora och små bokstäver i sökningen.  
Stor bokstav placeras före liten.  
Område innehåller kolumnhuvuden  
Om du har markerat den här rutan, ignoreras den första markerade tabellraden vid sorteringen.  
Inkludera format  
Om du inte har markerat den här rutan, är formateringarna av enskilda celler oförändrade efter en sortering.  
Detta är också fallet om innehållet i cellen ändras.  
Normalt är formateringar inte knutna till texten i en cell utan till själva cellen.  
Men om du har markerat den här rutan, binds formateringarna till texten i cellen och förflyttas till målpositionen vid en sortering.  
Sorteringsresultat till  
Om du har markerat den här rutan, placeras resultatet av en sortering i ett i förväg definierat tabellområde.  
Sorteringsresultat  
Om du har definierat ett tabellområde, kan du välja det här.  
Sorteringsresultat  
Här anger du cellområdet där sorteringsresultatet ska placeras.  
Användardefinierad sorteringsordning  
Om du markerar den här rutan, används en användardefinierad sorteringsordning.  
Om det tabellområde som ska sorteras innehåller begrepp som finns på den valda sorteringslistan, sorteras dessa med högsta prioritet och placeras alltså framför bokstaven A.  
Dessa begrepp sorteras i enlighet med sina förekomster i listan.  
Om du t.ex. har lagt in orden "januari, februari, februari januari" huller om buller i en tabellspalt och sorterar dem med en användardefinierad sorteringslista, får du resultatet "januari, februari, januari, februari ".  
Basen för den här sorteringsordningen är sorteringsalgoritmens arbetssätt.  
Den söker i den användardefinierade sorteringslistan efter "januari", hittar den termen och söker därefter inte från sorteringslistans början utan fortsätter på den plats där den senaste termen hittades.  
Användardefinierad sorteringsordning  
I den här listrutan väljer du en av de användardefinierade sorteringsordningarna som definierats under Verktyg - Alternativ - Tabelldokument...... - Sorteringslistor.  
Språk  
Språk  
Välj vilket språk som ska styra sorteringen.  
Alternativ  
Här väljer du ett alternativ för det valda språket.  
Riktning  
Uppifrån och ned (sortera rader)  
Om du väljer det här alternativet, sorteras alla rader i de markerade kolumnerna i det valda området.  
Från vänster till höger (sortera kolumner)  
Om du väljer det här alternativet, sorteras alla kolumner i de markerade raderna i det valda området.  
Dataområde  
Här visas det område som du har markerat för sortering.  
Filter  
Den här undermenyn innehåller kommandon för filtrering av data.  
Om du har definierat ett databasområde märker %PRODUCTNAME det automatiskt när markören står i en cell i området.  
Om markören står utanför ett databasområde så skapas ett namnlöst databasområde som används när kommandot utförs.  
Följande alternativ är tillgängliga:  
Standardfilter...  
Specialfilter...  
AutoFilter  
Med hjälp av AutoFilter kan du välja vissa värden från en datalista eller databas, som ska visas på kalkylarket.  
I listrutorna kan du välja vilka celler som ska filtreras ut.  
Välj posten -Standard - så öppnas dialogrutan Standardfilter.  
Där kan du ange ytterligare filtervillkor.  
Välj posten Top 10 om du bara vill visa de tio högsta värdena och dölja de övriga.  
Fler  
Om du klickar på den här kommandoknappen visas ett område där du kan välja bland olika funktioner för definition av filter.  
Alternativ  
Det här området innehåller olika inställningar.  
Versalkänslig  
Om den här rutan är markerad, gör programmet skillnad på stor och liten bokstav när filtret används på en lista.  
Område innehåller kolumnhuvuden  
Om den här rutan är markerad tas hänsyn till kolumnhuvudena på tabellens första rad.  
Skriv resultat till  
Om den här rutan är markerad kan du definiera ett utmatningsområde för resultatet av filteranvändningen.  
Du kan välja ett namngivet område i den enradiga listrutan.  
Du kan också markera ett område direkt på tabellarket som ska användas som utmatningsområde för filtreringsresultatet.  
AutoFilter-listrutorna visas då bara i det nya utmatningsområdet.  
Reguljärt uttryck  
Markera den här rutan om du vill använda platshållare vid filtreringen. %PRODUCTNAME stöder följande platshållare:  
Tecken  
Funktion / användning  
.  
Om du skriver "J.nsson" hittas "Jansson", "Jönsson "eller "Jonsson".  
^Peter  
Ordet hittas enbart om det står i början av ett stycke.  
Peter$  
Ordet hittas enbart om det står i slutet av ett stycke.  
*  
Med "Peter .*hemma" hittas t ex "Peter är hemma "och "Peter bor hemma".  
+  
Med "AX .+4" hittas "AX 4", men inte "AX4 "  
\t  
Hittar ett tabbtecken.  
()  
Med "(Peter har) _BAR_ (Peter får)" hittas både "Peter har "och "Peter får" i en sökning.  
\>  
Med "sol\>" hittas "vårsol "men inte "solsken".  
\<  
Med "\sol>" hittas "solsken "men inte "vårsol".  
Om de reguljära uttrycken är aktiverade, gäller de både för jämförelsen EQUAL (=) och för NOT EQUAL (<>).  
Detsamma gäller för funktioner som alltid arbetar med reguljära uttryck när det gäller strängar.  
DANTALV, DHÄMTA, PASSA, ANTAL.OM, SUMMA.OM, LETAUPP, LETARAD och LETAKOLUMN.  
Unika  
Den här funktionen utesluter dubbletter i utmatningsområdet efter en filtrering.  
Om samma resultat har filtrerats ut flera gånger reduceras alltså utmatningen till en (1) post.  
Behåll filterkriterier  
Om du markerar rutan Skriv resultatet till och anger ett målområde kan du med den här kryssrutan bestämma att målområdet ska förbli kopplat med källområdet.  
Källområdet måste redan vara definierat som dataområde under Data - Definiera område.  
Det på detta sätt definierade filtret kan du använda gång på gång via Data Uppdatera område.  
Markören måste då stå i källområdet.  
Dataområde  
Här anges det dataområde i tabellen på vilket filtret används i form av en referens.  
Om Du arbetar med ett känt område visas även dess namn här.  
Specialfilter  
I den här dialogrutan definierar du ett specialfilter.  
I ett specialfilter kan du kombinera upp till åtta olika filterkriterier.  
Filterkriterier finns i  
I listrutan väljer du områdesnamnet för det tabellområde, där det erforderliga filterkriteriet anges.  
Om du inte har gett det berörda området något namn så anger du området som innehåller filterkriteriet direkt i fältet till höger, eller markerar det aktuella området medan dialogrutan är öppen.  
Fler>>  
Ta bort filter  
Filtren i det markerade tabellområdet tas bort.  
Placera markören i det filtrerade cellområdet.  
Välj kommandot Ta bort filter.  
Samtliga filter som definierats gemensamt tas bort.  
Dölj AutoFilter  
Kommandoknapparna som du har definierat för AutoFilter för ett tabellområde visas inte längre.  
Detta påverkar inte AutoFiltrets funktion att dölja vissa rader.  
Delresultat  
I den här dialogrutan definierar du inställningar för automatisk beräkning av delresultat.  
Delresultat kan vara delsummor eller resultat av andra matematiska funktioner, som beräknas automatiskt i en tabell när ett värde i en viss kolumn i tabellen ändras.  
Om du har definierat ett databasområde märker %PRODUCTNAME det automatiskt om markören står i en cell i området.  
Om markören står utanför ett databasområde så skapas ett namnlöst databasområde som används när kommandot utförs.  
Då kan Du använda en delresultatfunktion för automatisk summering av omsättningen i de berörda postnummerområdena.  
Radera  
Med den här kommandoknappen raderar Du delresultatrader i ett markerat område.  
Grupp 1, 2, 3  
Här definierar du inställningarna för en av de tre delresultatsgrupperna.  
Alla delresultatflikar har samma struktur.  
Om du vill infoga delresultat för en tabell gör du på följande sätt:  
Markera först tabellen eller tabellområdet för vilket delresultat ska beräknas.  
I listrutan Gruppera efter väljer du sedan den kolumn där en värdeförändring automatiskt ska leda till en beräkning av ett delresultat.  
I rutorna i området Beräkna delresultat för väljer du en eller flera kolumner för vilka delresultaten ska beräknas med en funktion som du väljer i listrutan Beräkningsregler.  
Gruppera efter  
I den här listrutan väljer du den kolumn som ska styra beräkningsprocessen för delresultat.  
Om innehållet ändras från en rad till nästa inom den kolumn som Du anger här, utlöses beräkningen av ett delresultat automatiskt.  
Beräkna delresultat för  
I den här listrutan väljer du de markerade kolumner i tabellen vars cellinnehåll ska omfattas av beräkningen.  
Beräkningsregler  
I den här listrutan väljer fu den matematiska funktion som ska användas för beräkningen av delresultaten.  
Alternativ  
Här kan du göra några inställningar för hur delresultat beräknas och presenteras.  
Sidbrytning för varje grupp  
Om du markerar den här rutan påbörjas en ny sida efter varje delresultat.  
Versalkänslig  
Om du väljer det här alternativet leder även ändringar av stor och liten bokstav till att ett nytt delresultat skapas.  
Sortera området efter grupper först  
Om Du markerar den här kryssrutan sorteras det område som Du har angett på gruppflikarna under Gruppera efter enligt de angivna kolumnerna.  
Sortera  
I detta område anger Du alternativ för sorteringen av grupper.  
Inkludera format  
Om Du markerar denna kryssruta, tas även hänsyn till formateringar vid sorteringen.  
Användardefinierad sorteringsordning  
Om Du markerar den här kryssrutan, används en användardefinierad sorteringsföljd som Du har definierat på fliken Verktyg - Alternativ.. - Tabelldokument - Sorteringslistor och valt i listrutan.  
Stigande  
Om Du väljer detta alternativ sker sorteringen i stigande ordningsföljd, dvs från A till Ö och 0 till 9.  
Fallande  
Om detta alternativ valts sker sorteringen i fallande ordningsföljd, dvs från Ö till A och 9 till 0.  
Multipla operationer  
Med en multipel räkneoperation använder du samma formel på olika celler, men med olika värden som parametrar.  
För multipla operationer måste fältet Formler alltid vara ifyllt, medan bara ett av fälten Rad eller Kolumn måste innehålla en referens till den första cellen i respektive dataområde.  
Vid export till Microsoft Excel måste du tänka på att cellen med formeln bara får stå i vissa positioner i förhållande till dataområdet i Excel.  
Förinställningar  
Formler  
Här anger du en referens till cellerna, som innehåller de formler som den multipla räkneoperationen baseras på.  
Rad  
Här anger Du en referens till den cell, som ska användas som variabel parameter för de rader på vilka den multipla räkneoperationen ska användas.  
Kolumn  
Här anger Du en referens till den cell som ska användas som variabel parameter för de kolumner på vilka den multipla räkneoperationen ska användas.  
Konsolidera  
Med den här funktionen kan du sammanfatta data från flera fristående tabellområden.  
Med utgångspunkt från dessa områden räknar du sedan fram ett nytt område med hjälp av en matematisk funktion.  
Om du ska konsolidera flera tabellområden, som kan finnas i olika tabeller i tabelldokumentet, gör du så här:  
Först öppnar du dialogrutan för konsolidering.  
Med dialogrutan öppen markerar du de tabellområden som ska konsolideras och klickar på Lägg till efter varje område som du har markerat.  
Slutligen väljer du beräkningsregler i dialogrutan, och under Konsolidera efter väljer du det område där beräkningens resultat ska placeras.  
Därefter visas resultatet av konsolideringen.  
Beräkningsregler  
I den här listrutan väljer du den matematiska funktion som ska användas för beräkning av konsolideringen.  
Konsolideringsområden  
I det här fältet visas de dataområden som du redan har valt ut för konsolideringen.  
Källdataområde  
Om du redan har definierat områden med namn, kan du välja dem i listrutan och lägga till dem i listan Konsolideringsområden.  
I textfältet kan du skriva cellområden direkt och lägga till dem i listan Konsolideringsområden.  
Om du placerar markören i textfältet och sedan väljer tabellområden med musen, införs det markerade området i textfältet.  
Resultat vid  
Här väljer du den cell som ska utgöra resultattabellens övre vänstra hörn.  
Konsolideringstabellen visas sedan med början i denna cell.  
I listrutan kan du välja ett tidigare definierat område, skriva en celladress direkt eller markera en cell med musen, om markören står i textfältet till höger.  
Lägg till  
Om du klickar på den här kommandoknappen läggs den referens som finns under Källdataområde till på listan Konsolideringsområden.  
Fler>>  
Om du klickar på den här kommandoknappen, utvidgas dialogrutan Konsolidera med området Konsolidera efter och Alternativ.  
Konsolidera efter  
Konsolidera efter  
I det här området anger du om kolumnhuvuden eller radetiketter ska beaktas vid konsolideringen.  
Om någon av kryssrutorna är aktiverad, och om det förekommer olika kolumnhuvuden eller radetiketter i de enskilda tabellområdena, så genomförs separata konsolideringar för dessa kolumner eller rader.  
Om ingen av rutorna är markerad, konsoliderar programmet varje cell efter dess placering i tabellen utan att kontrollera om alla data verkligen passar ihop.  
Kolumnerna eller raderna i de områden som ska konsolideras måste alltså inte vara placerade i samma ordning.  
Så länge deras beteckningar överensstämmer kan de även vara placerade i någon annan ordning.  
Radetikett  
Om den här kryssrutan är aktiv så tas det hänsyn till radetiketter.  
Kolumnhuvuden  
Om den här kryssrutan är aktiv så tas det hänsyn till kolumnhuvuden.  
Alternativ  
Referensdata  
Om du aktiverar den här kryssrutan så länkas data i konsolideringsområdet med källdata.  
Om du ändrar data i källområdena, beräknas och anpassas resultaten i konsolideringsområdet automatiskt på nytt.  
Fler <<  
Klicka här om du vill stänga den utvidgade dialogrutan.  
Disposition  
Med kommandona på menyn Data - Disposition kan du utforma din tabell på ett överskådligt sätt.  
När du har grupperat tabellen kan du visa och dölja de enskilda områdena i tabellen genom att klicka på grupperingsikonerna i sidmarginalen.  
Gruppering...  
Upphäv gruppering...  
Dölj detalj  
Med detta kommando kan du dölja en dispositionsnivå i den grupperade tabellen  
Det innebär att en detalj i tabelldispositionen tillfälligt döljs, tills du visar den igen med kommandot Visa detalj.  
Visa detalj  
Med den här funktionen visar du dolda tabellområden igen.  
Då visas en detalj igen som du tidigare har dolt med kommandot Dölj detalj.  
Gruppering  
Här kan du gruppera ett markerat tabellområde.  
I dialogrutan definierar du grupperingen efter rader eller kolumner.  
Genom att klicka på de här ikonerna kan du visa eller dölja de grupperade områdena.  
Om du vill upphäva en gruppering använder du kommandot Upphäv gruppering.  
Aktivera för  
Här anger Du om grupperingen ska ske för rader eller kolumner.  
Rader  
Med det här alternativet samlas markerade rader till en grupp.  
Kolumner  
Med det här alternativet samlar Du markerade kolumner till en grupp.  
Upphäv gruppering  
Här tar du bort den understa nivån i den befintliga grupperingen som du infogat med kommandot Gruppering.  
Upphäv för  
Här väljer du vilken gruppering som ska upphävas.  
Rader  
Tar bort gruppegenskaper för tabellrader.  
Kolumner  
Tar bort gruppegenskaper för tabellkolumner.  
AutoDisposition  
Med det här kommandot väljer du en automatisk disposition av rader och / eller kolumner.  
Alla kolumner till vänster om en formel eller alla rader ovanför en formel sammanfogas, om formeln refererar till motsvarande celler.  
Titta t.ex. på följande tabell:  
januari  
februari  
mars  
1:a kvartalet  
april  
maj  
juni  
2:a kvartalet  
100  
120  
130  
350  
100  
100  
200  
400  
I cellerna för 1:a kvartalet och 2:a kvartalet står en summaformel för de tre cellerna till vänster om dem.  
AutoDispositionen delar in den här tabellen i de båda kvartalen.  
Ett streck visar dispositionsområdet.  
Streckets begynnelsepunkt är ett minustecken.  
Om du klickar på begynnelsepunkten sammanfattas dispositionsområdet.  
Minustecknet blir till ett plustecken.  
Om du klickar på det senare visas det dolda området igen.  
Du upphäver AutoDispositionen med Data - Disposition - Ta bort.  
Ta bort  
Med det här kommandot kan du upphäva grupperingar igen, vare sig de har gjorts manuellt eller med funktionen AutoDisposition.  
Datapilot  
Här visas en undermeny där du kan starta Datapiloten och uppdatera eller radera celler som beräknats av Datapiloten.  
Starta...  
Välj ut källa  
Datapiloten kan arrangera om dina tabelldata.  
Du kan med fördel använda datapiloten om du ska ordna data i en tvådimensionell tabell tre - eller flerdimensionellt.  
Den ger dig alltid tillgång till den datavy som du behöver för tillfället.  
Urval  
Här väljer Du en datakälla.  
Aktuell markering  
Data i ett cellområde i %PRODUCTNAME Calc-dokumentet används som källdata.  
När Du bekräftar Ditt val med OK öppnas dialogrutan Datapilot, där Du kan definiera layouten och hur Datapilotens resultat ska visas.  
Datakälla som är registrerad i %PRODUCTNAME  
Markera det här alternativet om Du vill använda en databastabell eller -sökning, som infogats i %PRODUCTNAME, som datakälla.  
De data som ska användas behöver inte importeras till %PRODUCTNAME Calc-dokumentetet.  
Om Du bekräftar det här alternativet med OK öppnas dialogrutan Välj ut datakälla, där Du kan definiera källan exakt.  
Extern källa / gränssnitt  
Om Du markerar det här alternativet kan Du använda en extern OLAP-server som källa.  
Om Du bekräftar Ditt val med OK öppnas dialogrutan Extern datakälla, där Du kan definiera OLAP-datakällan i detalj i rutorna "Service", "Källa", "Namn", "Användare" och "Lösenord ".  
Om Du bekräftar med OK öppnas dialogrutan Datapilot där Du kan definiera layouten och hur Datapilotens resultat ska visas.  
Information om OLAP hittar Du i den allmänna ordlistan för %PRODUCTNAME.  
Om Du skapar en Datapilot-tabell utifrån %PRODUCTNAME Calc-data läses talformaten in från första dataraden och läggs in på motsvarande sätt i Datapilot-tabellen.  
Välj ut datakälla  
I den här dialogrutan väljer Du en databas och den exakta datakällan.  
Urval  
Du använder området för att välja den datakälla som redan har angetts i %PRODUCTNAME %PRODUCTVERSION.  
Databas  
Listrutan visar alla anmälda och därmed valbara databaser.  
Datakälla  
Välj i denna lista en källa som hör till den angivna databasen.  
Typ  
Du väljer typ av källa i den här listrutan.  
Posterna Tabell, Sökning och SQL respektive SQL (Native) är tillgängliga.  
OK  
I den kan Du ange layouten och hur datapilotens resultat ska visas.  
Datapilot  
I den här dialogrutan definierar Du layouten och återgivning av datapilotens resultat.  
Layout  
Här bestämmer Du hur datapiloten ska bygga upp tabellen.  
Dra helt enkelt de visade fälten till layoutområdena "kolumn", "rad" och "data ".  
Du kan när som helst ändra ordningsföljden för de placerade fälten och flytta dem inom området med musen.  
Du kan även lägga tillbaka dem genom att dra dem från layoutområdet till de andra kommandoknapparna.  
Denna etikett innehåller förutom namnet även den formel som används för att skapa data i dataområdet.  
Genom att dubbelklicka på någon av kommandoknapparna i området Data öppnar Du dialogrutan Datafält.  
Där kan Du välja den använda matematiska formeln.  
Även om du dubbelklickar på något av fälten i området Rad eller Kolumn öppnas dialogrutan Datafält.  
Du kan sedan bestämma om %PRODUCTNAME ska räkna ut och visa delresultat eller inte.  
Fler>>  
Med den här kommandoknappen utökar Du dialogrutan med området Resultat.  
Om Du klickar en gång till på kommandoknappen stängs området igen.  
Resultat  
I detta alternativområde kan Du göra inställningar för datapilot-tabellens utdata.  
Utdata från  
Välj ett definierat område i listrutan.  
Markera sedan ett tabellområde med musen eller ange ett cellområde direkt i textfältet.  
Så kan Du även undvika att utvärderingstabellen skapas direkt under ursprungstabellen.  
Om inget utdataområde definieras, skapas datapilottabellen nedanför källområdet, oberoende av eventuella befintliga data.  
Ignorera tomma rader  
Om Du har markerat den här kryssrutan, ignoreras tomma rader i ursprungstabellen.  
Identifiera kategorier  
Om Du har markerat den här kryssrutan, läggs rader utan radetikett automatiskt till nästa högre kategori som har angetts genom en radetikett.  
Totalresultat kolumner  
Om det här fältet är aktiverat, visas totalresultatet av kolumnberäkningen.  
Totalresultat rader  
Om det här fältet är aktiverat, visas totalresultatet av radberäkningen.  
Filter  
I den här dialogrutan definierar Du logiska villkor för filtrering av data ur en tabell.  
Kriterier  
Här kan Du definiera ett standardfilter genom att ange typ av operator, fältets namn, ett logiskt villkor och ett värde respektive en kombination av argument.  
Operator  
För följande argument kan Du välja mellan de logiska operatorerna OCH och ELLER.  
Fältnamn  
Välj ur listrutan det fältnamn ur den aktuella tabellen som Du vill sätta in i argumentet.  
Här står kolumnnamnen om det inte finns några texter som fältnamn.  
Villkor  
Ur listrutan kan Du välja mellan flera relationsoperatorer med vars hjälp posterna i fälten Fältnamn och Värde länkas.  
Du kan välja mellan följande relationsoperatorer:  
Villkor:  
=  
lika med  
<  
mindre än  
>  
större än  
<=  
mindre än eller lika med  
>=  
större än eller lika med  
<>  
inte lika med  
Värde  
I den här listrutan listas alla de värden som är möjliga under Fältnamn.  
Välj ett värde som Du vill använda i filtret.  
Du kan även välja posterna -tom - eller -inte tom - om Du vill filtrera efter tomma eller inte tomma poster.  
Fler>>  
Alternativ  
Den här kommandoknappen öppnar ett område där Du kan välja bland olika alternativ för att definiera filtret.  
Alternativ  
I det här området hittar Du olika inställningsalternativ.  
Skiftlägeskänslig  
Om Du aktiverar det här alternativet, och filtret används på en lista, så görs det åtskillnad mellan versaler och gemener.  
Reguljärt uttryck  
Aktivera den här kryssrutan om Du vill arbeta med platshållare vid filtreringen. %PRODUCTNAME stöder för detta följande platshållare:  
Tecken  
Funktion / användning:  
.  
Om Du skriver "J.nsson" hittar Du "Jansson", "Jönsson "eller "Jonsson".  
^Peter  
Ordet hittas enbart om det står i början av ett stycke.  
Peter$  
Ordet hittas enbart om det står i slutet av ett stycke.  
*  
Med "Peter .*hemma" hittas t ex "Peter är hemma "och "Peter bor hemma".  
+  
Med "AX .+4" hittas "AX 4", men inte "AX4 "  
\t  
Hittar en tabulator.  
()  
Med "(Peter har) _BAR_ (Peter får)" hittas både "Peter har "och "Peter får" under en enda sökning.  
\>  
Med "sol\>" hittas "vårsol "men inte "solsken".  
\<  
Med "\sol>" hittas "solsken "men inte "vårsol".  
Om de reguljära uttrycken är aktiverade, gäller de både för jämförelsen EQUAL (=) och för NOT EQUAL (<>).  
Samma sak gäller för funktioner, som alltid arbetar med allmänna uttryck när det gäller strängar:  
DANTALV, DHÄMTA, PASSA, ANTAL.OM, SUMMA.OM, LETAUPP, LETARAD och LETAKOLUMN.  
Unika  
Denna funktion utesluter duplikat i utdataområdet efter användning av filtret.  
Om samma resultat har filtrerats ut flera gånger reduceras alltså utmatningen till en (1) post.  
Dataområde  
Här anges enligt skrivsättet för referenser dataområdet för den tabell på vilken filtret används.  
Om Du arbetar med ett känt område visas även dess namn här.  
Fler <<  
Med den här kommandoknappen döljer Du den utvidgade delen av dialogrutan.  
Datafält  
Dialogrutans utseende skiljer sig åt beroende på om du har öppnat dialogrutan genom att dubbelklicka på ett fält i området Data i Datapiloten eller genom att dubbelklicka på ett fält i områdena Rad eller Kolumn.  
Delresultat  
I det här området definierar du typen av delresultat.  
Inga  
Om du markerar det här alternativet beräknas inget delresultat.  
Detta är standardinställningen.  
Automatiskt  
Om du markerar det här alternativet beräknas delresultatet automatiskt.  
Användardefinierade  
Klicka på det här alternativet om du själv vill bestämma vilken typ av delresultat som ska beräknas.  
Sedan kan du välja typ av delresultat i listrutan i området Delresultat.  
Funktion  
Här kan du definiera vilken typ av delresultat som ska beräknas genom att klicka på posterna.  
Poster från det här fältet kan bara väljas om du har markerat alternativet Användardefinierade resp. om du har öppnat den här dialogrutan genom att dubbelklicka på ett fält i området Data i datapiloten.  
Visa objekt utan data  
Med den här rutan kan du ställa in om det ska infogas tomma rader resp. kolumner i utdatatabellen för de element i datakällan som inte innehåller några data.  
Namn:  
Detta är namnet på den kommandoknapp som du har dragit till något av områdena Kolumn, Rad eller Data.  
Uppdatera  
Med det här menykommandot uppdaterar du tabeller som du har skapat med Datapiloten.  
Detta kan vara nödvändigt om t.ex. utgångsdata har ändrats.  
Radera  
Med detta kommando raderar du datapilottabellen.  
Då raderas tabellen där cellmarkören befinner sig.  
Uppdatera område  
Här uppdaterar du data i tabellen om de har infogats från en extern databas.  
Detta innebär att ändringarna som du har gjort av dessa data i tabellen skrivs över, och att data övertas från en extern databas som eventuellt kan ha ändrats.  
Validitet  
I den här dialogrutan kan du definiera olika validitetskriterier för ett markerat tabellområde.  
Kriterier  
Här bestämmer du vilka värden som ska tillåtas för validitetskriterierna.  
Välj validitetens randvillkor för de markerade cellerna.  
Här kan du, med hjälp av alla inmatningsfält tillsammans, t.ex. definiera kriterier av typen: "Tal mellan 1 och 10" eller "Texter som inte är längre än 20 tecken ".  
Tillåt  
I den här listrutan väljer du vilken typ av villkor du ställer för cellernas data.  
Beroende på vilket villkor du har valt kan övriga alternativ i dialogrutan ändras.  
Du kan välja bland följande villkor:  
Villkor  
Effekt  
Varje värde  
Ingen begränsning  
Heltal  
Bara heltal som motsvarar villkoret.  
Decimal  
Alla tal som motsvarar villkoret.  
Datum  
Alla tal som motsvarar villkoret.  
De registrerade värdena formateras på motsvarande sätt när du öppnar dialogrutan nästa gång.  
Tid  
Alla tal som motsvarar villkoret.  
De registrerade värdena formateras på motsvarande sätt när du öppnar dialogrutan nästa gång.  
Textlängd  
Inmatningar vars längd motsvarar villkoret.  
Tillåt tomma celler  
Om du markerar den här rutan, så är även tomma celler tillåtna i området med de markerade cellerna.  
I annat fall måste varje cell innehålla ett värde.  
Data  
I den här listrutan väljer du typ av villkor.  
I övriga fall visas ett inmatningsfält som heter Värde, Minimum eller Maximum.  
Värde  
Här anger du värdet som dessa data måste motsvara enligt villkoret.  
Här anger du värdet som dessa data måste motsvara enligt villkoret.  
Om du t.ex. har valt "mellan" eller "inte mellan "under Data, matar du in minimivärdet här.  
Minimum  
Här anger du ett minimivärde.  
Maximum  
Här anger du ett maximivärde.  
Inmatningshjälp  
Här skapar du inmatningshjälp som du sedan har tillgång till vid markering av en cell.  
Erbjud inmatningshjälp vid markering av en cell  
Om du markerar det här fältet, så kommer den hjälp som du skriver in i området Innehåll att visas i dokumentet så snart du markerar cellen.  
Om du har skrivit in text i området Innehåll i dialogrutan och sedan avmarkerar det här fältet, så går den inskrivna texten förlorad.  
Innehåll  
Här definierar du innehållet i inmatningshjälpen.  
Rubrik  
Här anger du rubriken som ska visas som överskrift i fetstil i inmatningshjälpen.  
Inmatningshjälp  
Skriv in texten som ska visas under rubriken i området Inmatningshjälp.  
Infoga radbrytningar för hand på långa rader genom att trycka på Retur.  
Felmeddelande  
Här bestämmer du vilket felmeddelande som ska visas när ogiltiga värden matas in.  
Dessutom kan du bestämma att det ska startas ett makro i samband med ett felmeddelande.  
Visa felmeddelande när ogiltiga värden matas in  
Om du markerar det här fältet och ogiltiga värden matas in, så visas en text som du har definierat.  
I annat fall visas en standardtext som talar om att inmatningen är ogiltig.  
I båda fallen förkastas den ogiltiga inmatningen och cellens tidigare värde bibehålls om du väljer åtgärden "Stopp".  
Samma sak gäller för åtgärderna "Varning" och "Information "om du stänger varnings - eller informationsdialogrutan med Avbryt.  
Om du inte stänger dialogrutan med Avbryt utan med OK, så bibehålls det ogiltiga värdet.  
Innehåll  
Här definierar du felmeddelandets text eller en åtgärd.  
Åtgärd  
Välj antingen den typ av dialogruta som ska visas vid en felaktig inmatning, eller "Makro" om ett tidigare skrivet makro ska utföras vid felinmatning. (Se exempelmakro i slutet av filen).  
Åtgärden "Stopp" visar en dialogruta som bara kan stängas med OK.  
Den ogiltiga inmatningen förkastas.  
Åtgärderna "Varning" och "Information "visar en dialogruta som kan stängas med OK eller Avbryt.  
Om dialogrutan stängs med OK förkastas inte den ogitliga inmatningen.  
Genomsök...  
Om du klickar på den här kommandoknappen öppnas dialogrutan Makro där du kan välja ut ett makro som ska utföras vid ett felmeddelande.  
Rubrik  
Här anger du antingen namnet på ett makro som ska utföras vid felaktig inmatning eller rubriken på den dialogruta som ska visas.  
Felmeddelande  
Här skriver du in texten som ska stå i dialogrutan som visas vid felaktig inmatning.  
Exempelmakro:  
Function ExampleValidity( CellValue as String, TableCell as String)  
Dim msg as string  
msg = "Ogiltigt värde:" & "'"& CellValue &"'"  
msg = msg & "i tabell:" & "'"& TableCell &"'"  
MsgBox msg ,16 ," Felmeddelande "  
End Function  
Talformat: valuta  
Med den här ikonen visar du cellinnehållet i valutaformat.  
Talformat: valuta  
Se även Format - Cell - Tal angående formatering av cellinnehåll.  
Talformat: procent  
Med den här ikonen visar du cellinnehållet i procentformat.  
Talformat: procent  
Se även Format - Cell - Tal angående formatering av cellinnehåll.  
Du kan använda procenttecknet när du gör beräkningar med procenttal:  
1% motsvarar 0,01  
1 + 16% motsvarar 116% eller 1,16  
1%% motsvarar 0,0001  
Talformat: standard  
Med den här ikonen visar du cellinnehållet i standard-talformat.  
Talformat: standard  
Se även Format - Cell - Tal angående formatering av cellinnehåll.  
Talformat: lägg till decimal  
Med den här ikonen lägger du till en decimal i visningen av en eller flera markerade celler vid ett talformat.  
Talformat: lägg till decimal  
Talformat: radera decimal  
Med den här ikonen tar du bort den sista decimalen i visningen av en eller flera markerade celler vid ett talformat.  
Visningen uppdateras och avrundas till det minskade antalet decimaler.  
Talformat: radera decimal  
Tabellområde  
I tabellområdet visas adressen för cellen där cellmarkören står eller, om ett enkelt område är markerat, cellreferensen till området.  
Om du har markerat ett område som har ett namn, visas områdets namn här.  
När du skriver in en formel visas en lista över de tio senast använda funktionerna i den här listrutan.  
Du kan överföra en av de här funktionerna till inmatningsraden på formellisten genom att klicka på den.  
Programmet registrerar såväl inmatning med hjälp av Funktionsautopiloten som direkt inmatning.  
Men vid direkt inmatning registreras bara funktioner som inte står inom parentes, t.ex. som parametrar för andra funktioner.  
Tabellområdesfält  
Du kan skriva in en referens direkt.  
Om referensen gäller för en enskild cell (t.ex. F1) så placeras cellmarkören direkt på den och vyn ställs in så att cellen visas.  
Om du anger en områdesreferens (t.ex. enligt mönstret A1:C4) så markeras området och visas.  
Summa  
Klicka sedan på ikonen.  
Summafunktion  
%PRODUCTNAME känner igen ett cellområde, förutsatt att cellerna redan innehåller data.  
Sammanhängande dataområden summeras uppåt (kolumn) eller åt vänster (rad).  
Om det redan finns flera summafunktioner i kolumnen / raden kan de sammanfogas till totalsummor.  
Klicka på ikonen Överta om du vill överföra summaformeln på det sätt som den visas på inmatningsraden.  
Ikonen Summa visas bara när du inte har aktiverat inmatningsraden.  
Funktion  
Genom att klicka på den här ikonen anger du att du vill skriva in en formel.  
Placera cellmarkören i cellen där du vill infoga formeln.  
Klicka på den här ikonen på formellisten.  
Skriv in formeln i formellisten eller markera den eller de celler som ska ingå som cellreferens i formeln.  
Du kan växla fritt mellan att mata in via tangentbordet eller att markera celler med musen, beroende på vad som krävs för formeln.  
Den här ikonen är bara synlig om inmatningsraden inte är aktiverad.  
Funktion  
Inmatningsrad  
I den här delen av formellisten bygger du upp en formel.  
Du kan skriva in siffror eller text direkt som sedan infogas i cellen, eller själv skapa en formel med hjälp av Funktionsautopiloten.  
Inmatningsrad  
Ignorera  
Med det här kommandot ignorerar du ändringar i cellinnehållet.  
Det ursprungliga innehållet visas sedan på nytt i formelfältet.  
Ignorera cellinnehåll  
Överta  
Med det här kommandot överför du det aktuella innehållet från formelfältet till arbetsområdet.  
Detta infogas i den tabellcell som redigeras för tillfället.  
Klicka på den här ikonen när du vill avsluta redigeringen av tabellcellen.  
Överta  
Temaurval  
I dialogen Temaurval kan du byta ut vissa cellformatmallar.  
Cellformatmallarna som du kan byta ut är användarformatmallar (stilar) med fast angivna namn, som bl.a. bestämmer cellernas teckensnitt, inramning och bakgrundsfärg.  
Dialogrutan öppnas när du klickar på ikonen Temaurval på verktygslisten i ett %PRODUCTNAME Calc-dokument.  
Temaurval  
Klicka på en post i den stora listrutan.  
Resultatet visas omedelbart i den aktuella tabellen.  
Om du vill överta resultatet klickar Du på OK.  
Position i dokument  
Här visas numret för den aktuella tabellen och det totala antalet tabeller i dokumentet.  
Visningen sker enligt mönstret Tabell X / Y.  
X står för tabellens nummer i det aktuella dokumentet enligt tabellflikarnas ordningsföljd, från vänster till höger i nedre kanten av fönstret.  
Y står för det totala antalet tabeller i det aktuella dokumentet.  
Standardformel, datum / klockslag, felmeddelande  
I fältet längst till höger på statuslisten visas aktuell information om dokumentet.  
I normala fall visas standardformeln Summa här.  
Standardformeln Summa visar alltid summan av de markerade cellerna.  
Om ett fel har uppstått i den aktuella cellen visas felkoderna i klartext när cellen är markerad.  
På snabbmenyn för det här fältet på statuslisten kan du välja en annan standardformel.  
De tillgängliga alternativen är Medelvärde, Antal värden (ANTALV), Antal tal (ANTAL), Maximum, Minimum eller Inga.  
Om du väljer det sista alternativet visas datum och klockslag.  
Om du markerar hela rader eller kolumner med många tal så kanske det tar för lång tid att beräkna summan eller en annan funktion och visa resultatet på statuslisten.  
Då kan du välja alternativet Inga.  
Förstora skala  
Varje gång du klickar på den här ikonen förstoras förhandsgranskningen ett steg.  
Den aktuella skalan visas i skalafältet på statuslisten.  
Största skalan som kan användas är 400%.  
Förstora skala  
Minska skala  
Varje gång du klickar på den här ikonen förminskas förhandsgranskningen ett steg.  
Den aktuella skalan visas i skalafältet på statuslisten.  
Den minsta skalan som kan användas är 20%.  
Minska skala  
Infoga  
Med den här ikonen öppnar du en utrullningslist med funktioner för infogning av grafik och specialtecken.  
Ikon på verktygslisten:  
Infoga  
När du för första gången har valt en funktion på utrullningslisten, visas alltid ikonen för den senast infogade funktionen på utrullningslisten.  
Om du drar bort den från verktygslisten, får du tillbaka listen med dess olika funktioner.  
Du kan välja följande funktioner:  
Infoga grafik  
Infoga specialtecken  
Infoga celler  
Med den här ikonen öppnar du en utrullningslist med funktioner för infogning av celler, rader och kolumner.  
Ikon på verktygslisten:  
När du för första gången har valt en funktion på utrullningslisten, visas alltid ikonen för den senast infogade funktionen på utrullningslisten.  
Om du drar bort den från verktygslisten, får du tillbaka listen med dess olika funktioner.  
Du kan välja följande funktioner:  
Infoga celler, nedåt  
Infoga celler, till höger  
Infoga rader  
Infoga kolumner  
Kortkommandon för tabelldokument  
Här hittar du tangentkommandon som är specifika för tabelldokument.  
Dessutom gäller de allmänna tangentkombinationerna i %PRODUCTNAME.  
Du använder tangentkombinationen Alternativ Alt +Retur i tabelldokument för att fylla i ett markerat område med den aktuella cellens innehåll.  
Markera ett område i tabellen, ange ett värde eller en formel och avsluta med den här tangentkombinationen.  
Hela det markerade området fylls i.  
Om du använder tangentkombinationen Skift Kommando +Ctrl +Retur när du har markerat ett område och skrivit in ett värde eller en formel, definierar du ett matrisområde, där alla celler får innehållet som du har skrivit in.  
Ett matrisområde är skyddat mot ändringar av dess delar.  
Du kan använda tangenten Kommando Ctrl som funktionstangent när du markerar celler med musen och vill göra en delad markering.  
De celler som du markerar med musen när du håller ner Ctrl-tangenten utgör en delad markering.  
Om du vill redigera eller skriva ut flera tabeller i det aktuella dokumentet samtidigt kan du markera dem gemensamt:  
Håll ner Kommando Ctrl -tangenten och klicka på tabellflikarna nedtill i dokumentfönstret.  
En ljus tabellflik visar att tabellen är markerad och en grå tabellflik att tabellen inte är markerad.  
På snabbmenyn finns även ett kommando för att markera alla tabeller.  
Om du håller ner skifttangenten och klickar på fliken för den aktuella tabellen markeras bara den aktuella tabellen.  
Med tangentkombinationen Kommando Ctrl +Retur infogar du en manuell radbrytning direkt i en cell (inte på inmatningsraden).  
Då bryts texten automatiskt i den högra kolumnkanten.  
Där väljer du vilket innehåll du vill radera i cellen.  
Med backstegstangenten (ovanför returtangenten) raderar du innehållet i cellen utan dialogruta.  
Navigera i tabelldokument  
Tangentkombination  
Effekt  
Kommando Ctrl +Home  
Placerar markören i cell A1  
Kommando Ctrl +End  
Placerar markören i den sista cellen som innehåller data i det aktuella tabelldokumentet.  
Om den sista raden med data är rad 10 och den sista kolumnen med värden är kolumn F, placeras markören i cell F10.  
Home  
Placerar markören i kolumn A på den aktuella raden.  
End  
Placerar markören i den sista kolumnen med data på den aktuella raden.  
Kommando Ctrl +x  
* är multiplikationstecknet på den numeriska delen av tangentbordet  
Markerar hela blocket där markören står.  
Ett block är ett sammanhängande område av celler som är fyllt med data.  
Retur i ett markerat block  
Placerar markören i nästa cell inne i ett block.  
Markörens riktning kan ställas in under Verktyg - Alternativ - Tabelldokument - Allmänt.  
Kommando Ctrl +Vänsterpil  
Hopp till den vänstra kolumnen i det aktuella blocket eller hopp till föregående block.  
Om det inte finns något block, hopp till den första kolumnen, A.  
Kommando Ctrl +Högerpil  
Hopp till den högra kolumnen i det aktuella blocket eller hopp till nästa block.  
Om det inte finns något block, hopp till den sista kolumnen, IV.  
Kommando Ctrl +Uppåtpil  
Hopp till den översta raden i det aktuella blocket eller hopp till föregående block.  
Om det inte finns något block, hopp till den första raden, 1.  
Kommando Ctrl +Nedåtpil  
Hopp till den understa raden i det aktuella blocket eller hopp till nästa block.  
Om det inte finns något block, hopp till den sista raden, 32000.  
Kommando Ctrl +Page Up  
Hopp till föregående tabellark  
I förhandsgranskningen: hopp till föregående utskriftssida.  
Kommando Ctrl +Page Down  
Hopp till nästa tabellark  
I förhandsgranskningen: hopp till nästa utskriftssida.  
Alternativ Alt +Page Up  
Rullar en bildskärmssida åt vänster  
Alternativ Alt +Page Down  
Rullar en bildskärmssida åt höger  
Tabelldokumentsfunktioner med funktionstangenterna  
Tangentkombination  
Effekt  
F2  
Växla till redigeringsläge  
Kommando Ctrl +F2  
Öppna Funktionsautopiloten  
F3  
Infoga namn  
Kommando Ctrl +F3  
Öppna dialogrutan Definiera namn  
F4  
Visa / dölj aktuell databas  
Skift+F4  
Växla mellan relativa / absoluta referenser i inmatningsfält (A1, $A$1, $A1, A$1)  
F5  
Navigator  
Skift+F5  
Visa spår till efterträdaren  
Kommando Ctrl +F5  
Visa spår till föregångaren  
F7  
Öppna rättstavningskontrollen  
Kommando Ctrl  
Öppna synonymordlistan  
F8  
Kompletteringsläge på / av  
Skift+F8  
Utökningsläge på / av  
Kommando Ctrl +F8  
Framhäv värden  
F9  
Beräkna på nytt  
Kommando Ctrl +F9  
Uppdatera diagram  
F11  
Stylist  
Skift+F11  
Skapa mall  
Skift + Kommando Ctrl +F11  
Uppdatera mall  
F12  
Gruppering på  
Kommando Ctrl +F12  
Gruppering av  
Formatering av tabelldokument med kortkommandon  
Följande cellformat kan ställas in direkt med kortkommandon:  
Tangentkombination  
Effekt  
Kommando Ctrl +Skift+1 (inte på den numeriska delen av tangentbordet)  
Två decimaler, tusentalsavgränsare  
Kommando Ctrl +Skift+2 (inte på den numeriska delen av tangentbordet)  
Standardformat för exponent  
Kommando Ctrl +Skift+3 (inte på den numeriska delen av tangentbordet)  
Standardformat för datum  
Kommando Ctrl +Skift+4 (inte på den numeriska delen av tangentbordet)  
Standardformat för valuta  
Kommando Ctrl +Skift+5 (inte på den numeriska delen av tangentbordet)  
Standardformat för procent (2 decimaler)  
Kommando Ctrl +Skift+6 (inte på den numeriska delen av tangentbordet)  
Standardformat  
Kommando Ctrl +*  
* är multiplikationstecknet på den numeriska delen av tangentbordet  
Markerar det aktuella området  
Alternativ Alt +Nedåtpil  
Den aktuella raden blir högre  
Alternativ Alt +Uppåtpil  
Den aktuella raden blir lägre  
Alternativ Alt +Högerpil  
Den aktuella kolumnen blir bredare  
Alternativ Alt +Vänsterpil  
Den aktuella kolumnen blir smalare  
Alternativ Alt +Skift+Piltangent  
Ställer in optimal kolumnbredd eller radhöjd efter innehållet i den aktuella cellen.  
Felkoder i %PRODUCTNAME Calc?  
Här lär du dig vad felkoderna i %PRODUCTNAME Calc betyder.  
Här får du förutom felmeddelandet även själva feltexten och en kort förklaring av felet.  
Felkoden visas tillsammans med hänvisningen Err:.  
Om den cell som innehåller felet är aktiv, så visas feltexten i statuslisten.  
Felkod  
Feltext  
Förklaring  
501  
Ogiltigt tecken  
Ett tecken som är ogiltigt i detta sammanhang, t ex =1Eq i stället för =1E2  
502  
Ogiltigt argument  
En funktions argument har ett ogiltigt värde, t ex ett negativt tal vid funktionen ROT()  
503  
Ogiltig flyttalsoperation  
T ex division med 0 eller andra beräkningar som orsakar ett spill där den definierade värdemängden överskrids  
504  
Fel i parameterlistan  
Någon parameter i en funktion är av ogiltig typ, t ex text i stället för tal, eller områdesreferens i stället för enskild cellreferens  
505  
Internt syntaxfel  
Används inte  
506  
Ogiltigt semikolon  
Används inte  
507  
Felplacerade parenteser  
Används inte  
508  
Felplacerade parenteser  
T ex avslutande parentes utan tillhörande inledande parentes, eller att avslutande parentes saknas inuti formeln (saknad avslutande parentes i slutet av formeln tillfogas automatiskt)  
509  
Operator saknas  
T ex =2( 3+4) * mellan 2 och (bortglömd operator  
510  
Variabel saknas  
Två operatorer, varav den andra inte är någon enställig operator, följer direkt efter varandra, t ex =1+*2  
511  
Variabel saknas  
Funktionen behöver fler variabler än vad som har angetts, t ex OCH() och ELLER() utan parameter  
512  
Formel för lång  
Kompilator: som redan namnet skvallrar om... syftar till det interna antalet symboler (max 512).  
Detta antal har inget att göra med den inmatade formelns stränglängd utan avser antalet operatorer, variabler, parenteser etc.  
Tolk: formler som skapar för många matriser på en gång (max 150), även Basic-funktioner som får för stor matris som parameter (max 0xFFFE, alltså 65534 byte)  
513  
Sträng för lång  
Kompilator: en identifierare i formeln är större än 64KB.  
Tolk: ett resultat till en strängoperation är större än 64KB  
514  
Internt spill  
Sorteringsoperationer med för många numeriska data (max 100000) eller spill i räknestacken.  
515  
Internt syntaxfel  
Används inte  
516  
Internt syntaxfel  
En matris förväntas på räknestacken, men finns inte där  
517  
Internt syntaxfel  
Okänd OpCode, t ex ett dokument med en ny funktion som laddats i en gammal version som ännu inte har denna funktion  
518  
Internt syntaxfel  
En variabel som ska flyttas ut från räknestacken finns inte  
519  
inget resultat (I cellen står inte Err:519 utan #VÄRDE!)  
En funktion har inte kunnat leverera ett värde som motsvarar definitionen, eller en cell som formeln refererar till innehåller text i stället för ett tal som behövs  
520  
Internt syntaxfel  
Kompilatorn har skapat kod som är okänd för den själv  
521  
Internt syntaxfel  
Inget resultat på räknestacken  
522  
Cirkelreferens  
En formel hänvisar direkt eller indirekt till sig själv och under Verktyg / Alternativ / Tabelldokument / Beräkna är iterationerna inte aktiverade  
523  
Beräkningssätt konvergerar inte  
En del (finans - )statistiska funktioner som måste närma sig ett visst värde, men som inte gör det, eller iterationer av cirkelreferenser som inte uppnår den minsta ändringen inom det inställda maximala antalet steg  
524  
Ogiltig referens (i cellen står inte Err:524 utan #REF!)  
Kompilator: ett kolumn - / radetikettnamn har inte kunnat lösas upp.  
Tolk: i formeln refereras till en cell vars kolumn, rad eller tabell har raderats, eller som skulle ligga utanför  
525  
Ogiltigt namn (i cellen står inte Err:525 utan #NAMN?)  
En identifierare kunde inte utvärderas( exempel: ingen giltig referens, inget giltigt områdesnamn, ingen kolumn - / radetikett, inget makro, fel decimaltecken, add-in hittades inte).  
526  
Internt syntaxfel  
föråldrad, används inte längre, men skulle dock kunna komma från gamla dokument om en formels resultat är ett område  
527  
Internt spill  
Tolk: för djup kapsling av referenser (en cell refererar till en cell, som refererar till en cell, som refererar till en cell osv)  
Känna igen namn som adressering  
%PRODUCTNAME kan i stor utsträckning tilldela områden namn självständigt under förutsättning att du har angett rad - och kolumnetiketter.  
Se följande tabell:  
Den automatiska namnidentifieringen gör det möjligt att mata in formeln =SUMMA( juli) i cell B8 i vårt exempel.  
I cell C8 blir den till =SUMMA( augusti) och i D8 till =SUMMA(september).  
Den här hjälpen fungerar även i horisontell riktning:  
Mata till exempel in formeln =SUMMA( London) i cell E4.  
Eftersom det här namnet innehåller mellanslag, måste det omges med enkla citationstecken (apostrofer): =SUMMA('New York').  
Den automatiska identifieringen arbetar inte med formler.  
Du kan alltså inte mata in formeln =SUMMA( Summa) i cell E8 men däremot =SUMMA(B8:D8) eller =SUMMA(E3:E6).  
Den sistnämnda formeln sätts för övrigt även in om du placerar markören i cell E8 och helt enkelt klickar på summaikonen på formellisten.  
Funktionen är aktiverad som standard.  
Du kan deaktivera den under Verktyg - Alternativ... - Tabelldokument - Beräkna.  
Ta bort markeringen i fältet Sök kolumn - / radetiketter automatiskt.  
Om du vill ha mer kontroll över namnen definierar du dem själv med kommandot Infoga - Namn - Etiketter....  
För att namn skall identifieras automatiskt som beteckningar måste de bestå av alfanumeriska tecken och det första tecknet måste vara en bokstav.  
Om du även vill använda icke-alfanumeriska tecken, inklusive mellanslag, måste du skriva namnet med enkla citationstecken (').  
Om en apostrof förekommer i namnet, som t.ex. i jan '97, måste ett omvänt snedstreck stå framför det här tecknet (jan \'97).  
Denna typ av referens är inte kompatibel med tidigare versioner av %PRODUCTNAME.  
Adressering med namn  
En elegant lösning för att göra referenserna till celler och cellområden i formler mer läsbara är att ge områdena namn.  
Kalla t.ex. området A1:B2 för Start.  
Du kan sedan helt enkelt skriva "=SUMMA(Start)" i formeln. %PRODUCTNAME tilldelar de namngivna områdena korrekt även när du har infogat eller raderat rader och kolumner.  
Områdesnamn får inte innehålla mellanslag.  
Om du till exempel har utvecklat en formel för beräkning av mervärdesskatt, så är det säkert lättare att läsa om du skriver "= Belopp * Skattesats" i stället för till exempel "= A5 * B12 ".  
Här skulle du ha kallat cell A5 för "Belopp" och cell B12 för "Skattesats ".  
Mata in namnet på det första området och klicka på Lägg till.  
I dialogrutan kan du även definiera fler namn genom att först mata in namnet i textfältet och sedan markera cellerna som skall ha namnet i tabellerna.  
Använd även dialogrutan Definiera namn till att definiera formler eller delar av formler som du ofta använder med ett namn.  
Stäng dialogrutan med OK.  
Infoga tabell  
1.  
Peka med musen på tabellfliken i den undre fönsterkanten.  
2.  
Du ser kommandon för att redigera tabellerna.  
3.  
Dialogrutan Infoga tabell öppnas.  
4.  
Välj position och antal tabeller som ska infogas och klicka på OK.  
Dialogrutan Infoga tabell  
Fylla i celler automatiskt  
Om du markerar ett cellområde och sedan tar tag i den lilla rutan i områdets högra, nedre hörn med musen och drar ut den nedåt eller åt höger, fylls innehållet i de nya cellerna i automatiskt.  
Följden 1 2 blir till 1 2 3 4 osv., följden 1 3 blir till 1 3 5 7 osv., cellinnehållet "1 kvartalet" blir till 1 kvartalet 2 kvartalet 3 kvartalet o.s.v., cellinnehållet "avdelning 1 "blir till avdelning 1 avdelning 2 avdelning 3 osv.  
Tal ändras alltså men inte texter.  
De texter som finns i sorteringslistorna (meny Verktyg - Alternativ - Tabelldokument - Sorteringslistor) utgör ett undantag.  
Om du t.ex. börjar dra serien jan feb med musen, fylls serien i med förkortningar av månadsnamnen.  
Om värdena inte ska ändras automatiskt håller du ner Kommando Ctrl -tangenten medan du drar.  
Hur kan ett datumfält fortsätta automatiskt med nästa månad i en kolumn i ett tabelldokument?  
För in 01.01.00 i cell A1  
För in 01.02.00 i cell A2  
Markera båda fälten med musen (så att båda är markerade samtidigt).  
I cell A2 ser du en liten kvadrat i det högra undre hörnet av cellen.  
För muspekaren till den här kvadraten tills markören förvandlas till ett kors.  
Dra sedan musen neråt (så att flera fält i kolumnen markeras).  
Om du nu släpper musknappen fylls fälten i kolumnen med datum där respektive månad är angiven.  
Använda AutoFilter  
Funktionen AutoFilter skapar listor i kolumnerna, där du väljer vilka dataposter (rader) som ska visas.  
Markera ett tabellområde som ska filtreras.  
Välj Data - Filter - AutoFilter.  
Listrutorna visas i den första raden i det markerade området.  
Välj ett värde i en listruta.  
Bara de rader visas vars innehåll motsvarar filterkriterierna.  
De andra raderna döljs.  
Du kan se att rader är dolda på avbrottet i radnumren.  
Kolumnen som använts för filtreringen markeras med en annan färg på pilknappen.  
Om du väljer posten -alla - i AutoFilter-listrutan i en cell visas alla rader igen.  
Om du vill ta bort listrutorna markerar du alla celler som du markerade i steg 1 och väljer kommandot Data - Filter - AutoFilter igen.  
I %PRODUCTNAME Calc tar beräkningsfunktionen även med dolda celler.  
Summman av en hel kolumn summerar t.ex. även värdena i de dolda cellerna.  
Använd funktionen DELSUMMA om bara de celler som är synliga när du har använt ett filter ska tas med i beräkningen.  
Data - Filter - AutoFilter  
DELSUMMA  
Använda AutoFormat för tabell  
En snabb möjlighet att formatera en tabell eller ett cellområde finns i funktionen Format - AutoFormat.  
Markera först cellerna som skall formateras automatiskt, inklusive kolumn - och radhuvudena och eventuell summarad eller -kolumn.  
Minst 3x3 celler måste vara markerade innan den här menypunkten aktiveras.  
Sedan öppnar du dialogrutan AutoFormat.  
I förhandsvisningsområdet ser du ett exempel på hur respektive formatering som du väljer i fältet Format skulle se ut.  
Klicka på OK för att använda formateringen på det markerade området i tabellen.  
Om du inte ser färgändringar av cellinnehållet, är det möjligt att Framhäv värden är markerat under Verktyg - Alternativ - Tabelldokument - Vy - Visa eller på menyn Visa.  
I så fall används de förinställda färgerna.  
Du kan definiera dina egna formateringar som AutoFormat:  
Formatera en tabell som du vill  
Markera hela den formaterade tabellen, genom att t.ex. klicka på kommandoknappen utan text till vänster ovanför radhuvudena.  
Öppna dialogrutan AutoFormat och klicka där på Lägg till.  
Du definierar sedan ett namn för det nya formatet i en dialogruta.  
I framtiden kan du även använda det egna AutoFormatet som du har definierat till andra tabeller.  
Du kan skapa mycket tilltalande tabeller för automatisk formatering genom att välja en lämplig bakgrundsfärg för tabellcellerna.  
Här kan du välja vilka av det valda formatets egenskaper som skall undantas från den automatiska formateringen.  
Om du till exempel tar bort markeringen i fältet Teckensnitt, påverkas inte teckensnitt vid automatisk formatering med AutoFormat.  
Format - AutoFormat  
Stänga av automatiska ändringar  
%PRODUCTNAME Calc korrigerar ett antal skrivvanliga fel enligt förinställningen.  
Du kan ångra varje automatisk ändring direkt, t.ex. med Kommando Ctrl +Z.  
Här följer ställena i %PRODUCTNAME där du stänger av automatiska ändringar (och sätter på dem igen):  
Text eller tal kompletteras automatiskt  
När du gör en inmatning i en cell kan %PRODUCTNAME Calc automatiskt upprepa en inmatning som förekommer i samma kolumn.  
Den här funktionen kallas AutoInmatning.  
Du sätter på resp. stänger av AutoInmatning genom att sätta en bock resp. ta bort den framför kommandot Verktyg - Cellinnehåll - AutoInmatning.  
Citatationstecken ersätts med typografiska anföringstecken  
Öppna ett tabelldokument.  
Välj Verktyg - AutoKorrigering.  
Klicka på fliken Typografiska anföringstecken.  
Avmarkera Ersätt.  
Cellinnehåll börjar alltid med stor bokstav  
Öppna ett tabelldokument.  
Välj Verktyg - AutoKorrigering.  
Klicka på fliken Alternativ.  
Avmarkera Börja varje mening med stor bokstav.  
Ord ersätts med ett annat ord  
Öppna ett textdokument.  
Välj Verktyg - AutoKorrigering.  
Klicka på fliken Ersättning.  
Leta upp ordparet och radera det.  
Verktyg - Cellinnehåll - AutoInmatning  
Verktyg - AutoKorrigering  
Räkna med datum och tid  
I tabelldokument kan du inte bara se datum och tid (de övertas från systemtiden på din dator).  
Du kan också räkna med datum - och tidsangivelser.  
Om du vill få reda på hur gammal du är i sekunder eller timmar, så gör du på följande sätt:  
Öppna ett nytt tomt tabelldokument.  
Skriv in ditt födelsedatum i cell A1, till exempel 64-09-04.  
Mata in följande formel i A3: =NU( )-A1.  
Så fort du trycker på returtangenten eller klickar på kommandoknappen Överta (den gröna bocken) ser du resultatet som automatiskt är formaterat som datum.  
Eftersom du vill se differensen mellan två datumangivelser som antal dagar, måste du formatera cellen A3 som tal.  
Placera markören i cell A3 och formatera cellen som tal.  
För att göra det öppnar du snabbmenyn i cell A3 (tryck på högra musknappen) och väljer Formatera celler...  
Du ser dialogrutan Cellattribut med fliken Tal där kategorin Tal är förinställd.  
Formatet är "Standard" vilket bland annat innebär att resultatet av en beräkning med datumangivelser visas som datum.  
Om du vill framtvinga visning som tal sätter du talformatet till t.ex. "-1.234" och stänger dialogrutan med OK.  
I cell A3 ser du nu antalet dagar mellan dagens datum och det inmatade datumet.  
Mata även in de andra formlerna om du vill: =A3*24 för timmar i A4, =A4*60 för minuter i A5 och =A5*60 för sekunder i A6 och bekräfta inmatningen som beskrivet ovan.  
Du ser nu att tiden sedan din födelsedag har beräknats och förts in i de olika enheterna.  
Värdet i sekunder refererar till tidpunkten då du bekräftade din formel i cell A6 med t.ex. returtangenten.  
Det här värdet uppdateras inte trots att "nu" ständigt fortsätter.  
På menyn Verktyg finns visserligen kommandot Cellinnehåll - Automatisk beräkning som är aktiverat enligt standard, men den här automatiken påverkar inte funktionen NU: din dator skulle i så fall bara vara upptagen med att uppdatera tabellen.  
Men för skojs skull kan du trycka på funktionstangenten F9 upprepade gånger för att beräkna tabellen på nytt.  
Låt fingret vila på F9 och se hur tiden rinner iväg.  
Beräkna serier automatiskt  
Mata in ett tal i en cell.  
Dra det högra undre hörnet på cellen nedåt med musen.  
När du släpper musknappen fylls cellerna som du har markerat med tal.  
Det här talet ökas med 1 för varje cell.  
Om du har markerat två eller flera angränsande celler som innehåller olika tal och drar upp dem gemensamt, fortsätter ett eventuellt aritmetiskt mönster av talen om ett sådant går att känna igen.  
Ett exempel:  
Om talet 1 står i A1 och talet 3 i A2 så fortsätter serien med 5, 7, 9, 11 och så vidare när du kopierar båda cellerna gemensamt genom att dra neråt.  
Markera först området som du vill fylla i tabellen.  
I dialogrutan som du nu kan öppna med Redigera - Fyll - Serie, väljer du typ av seriestruktur.  
Välj till exempel 2 som startvärde, 2 som inkrement och den geometriska serien som serietyp.  
Då får du en lista över potenserna av 2.  
Som du ser i den här dialogrutan kan du också fylla i datum - och tidsserier.  
Om du till exempel behöver den första i alla månader på året som radhuvuden, gör du på följande sätt:  
Mata till exempel in "00-01-01" i en cell (utan citationstecknen).  
Markera den här cellen och de 11 angränsande cellerna under den.  
Välj Redigera - Fyll - Serie.  
I dialogrutan väljer du alternativen Datum och Månad.  
Klicka på OK.  
Du ser nu datumet för första dagen i varje månad.  
Sorteringslistor  
Beräkna tidsskillnad  
Om du vill beräkna tidsskillnader, t.ex. hur lång tid det är mellan klockslagen 23:30 och 01:10 samma natt, kan du använda följande formel:  
=( B2<A2 )+B2-A2  
Det senare klockslaget står då i B2 och det tidigare klockslaget i A2.  
1 timme och 40 minuter.  
Formeln använder sig av att en hel dag med sina 24 timmar har värdet 1, och att en timme uppgår till 1 / 24 av detta värde.  
Det logiska värdet inom parentes är 0 eller 1, motsvarande 0 eller 24 timmar.  
Formelns resultat matas automatiskt ut i tidsformat p.g.a. operandernas ordningsföljd.  
Räkna i tabeller  
Följande enkla procenträkningsexempel visar hur du kan räkna i ditt tabelldokument:  
1.  
Placera cellmarkören i cellen A3.  
2.  
Skriv in talet 150 och tryck på returtangenten.  
Cellmarkören växlar neråt till cell A4.  
3.  
Mata in talet 16 i cell A4.  
Tryck inte på returtangenten den här gången, utan på tabb-tangenten.  
Cellmarkören växlar åt höger till cellen bredvid, B4.  
4.  
I cell B4 matar du in följande:  
=A3 * A4 / 100 "  
Om du inleder en inmatning med ett likhetstecken, så visar du att du vill mata in en formel.  
Du ser formeln på inmatningsraden på formellisten.  
5.  
Tryck på returtangenten för att avsluta formeln.  
Resultatet av beräkningen, nämligen 16 procent av 150 ser du som innehåll i cell B4.  
6.  
Klicka i cell A3, mata in 200 och tryck på returtangenten.  
Du ser att resultatet av beräkningen har anpassats automatiskt.  
7.  
Klicka i cell B4 och sedan vid slutet av formeln på inmatningsraden på formellisten.  
En blinkande textinmatningsmarkör visar att du kan göra en ny inmatning.  
8.  
Tillfoga "+ A3" (utan citationstecken) vid formelns slut och tryck på returtangenten.  
I cell B4 ser du nu det nya beräknade värdet av formeln: de tidigare beräknade 16 procenten av värdet från A3 plus innehållet i A3.  
Bara kopiera synliga celler  
Nu vill du bara kopiera de celler som fortfarande är synliga till ett annat ställe.  
%PRODUCTNAME hanterar celler olika beroende på hur du har dolt cellerna och vad du vill göra med dem.  
Metod  
Resultat  
Celler har filtrerats bort med AutoFilter, standardfilter eller specialfilter.  
Du kopierar de synliga cellerna, t.ex. med kommandona Kopiera och Klistra in via urklippet eller med musknappen i mitten eller med dra-och-släpp samtidigt som du håller ner Ctrl-tangenten.  
Bara cellerna som fortfarande är synliga kopieras.  
Celler har filtrerats bort med AutoFilter, standardfilter eller specialfilter.  
Du flyttar de synliga cellerna, t.ex. med kommandona Klipp ut och Klistra in via urklippet eller med dra-och-släpp.  
Alla celler, även de dolda, flyttas.  
Celler har dolts manuellt med kommandot Dölj på snabbmenyn till radhuvudena eller kolumnhuvudena eller genom en disposition.  
Du kopierar eller flyttar de synliga cellerna.  
Alla celler, även de dolda, kopieras eller flyttas.  
Skydda celler mot ändringar  
I standardinställningen är cellskyddet aktiverat för alla celler.  
Men det får bara effekt om du skyddar tabellen eller dokumentet.  
1.  
Om det finns celler som du inte vill skydda, t.ex. där användaren ska göra inmatningar, markerar du de här cellerna och upphäver deras cellskydd.  
Om du sedan skyddar tabellen eller dokumentet är alla andra celler skyddade mot ändringar.  
2.  
Välj Format - Cell och klicka på Cellskydd.  
Kryssrutorna under den här fliken är tristate-fält, som kan anta tre lägen.  
Om rutan är tom, gäller funktionen inte för någon av de markerade cellerna.  
Om rutan är markerad med en svart bock på vit grund, gäller funktionen för alla markerade celler.  
Om bocken och grunden är gråa, gäller funktionen för minst en cell, men inte för alla.  
3.  
Välj de funktioner som ska gälla för de markerade cellerna.  
Skyddad innebär att cellens innehåll och dess formatering inte kan ändras.  
Dölj formel innebär att de använda formlerna inte är synliga och inte kan ändras.  
På detta sätt kan den som utvecklar tabellformatmallar skydda sitt arbete mot obehörig insyn.  
Dölj vid utskrift innebär att cellerna syns på bildskärmen, men inte på papper.  
4.  
Stäng dialogrutan med OK.  
5.  
Du aktiverar skyddet genom att välja Verktyg - Skydda dokument och sedan antingen Tabell eller Dokument.  
Då visas en dialogruta där du kan ange ett lösenord.  
Skyddet träder i kraft om du avslutar den här dialogrutan med OK, även om du inte anger något lösenord.  
Om du anger ett lösenord och sedan glömmer bort det, finns det ingen möjlighet att upphäva skyddet igen!  
Därför är det bäst att inte ange något lösenord om du bara vill skydda cellerna mot oavsiktliga ändringar - då kan skyddet upphävas igen när som helst.  
Cellreferens med dra-och-släpp  
Med hjälp av Navigator kan du skapa en referens till celler från ett tabelldokument i en annan tabell i samma dokument eller i ett annat dokument.  
Cellerna kan infogas som kopia, som länk eller som hyperlänk.  
Området som ska infogas måste definieras i ursprungsfilen som område med ett namn så att det kan infogas i målfilen.  
Öppna dokumentet där källcellerna finns.  
Källområdet ska vara definierat som område, du kan t.ex. markera cellerna och välja Infoga - Namn - Definiera.  
Om du definierar området först nu sparar du källdokumentet en gång till.  
Öppna dessutom tabellen, där du vill infoga ett objekt, som aktuell tabell.  
Välj källfilen i det undre kombinationsfältet i Navigator.  
I Navigator ser du nu objekten som finns i källfilen, bl.a. även de områden som har definierats där.  
Välj om du vill ha en referens i form av hyperlänk, länk eller kopia med ikonen Draläge i Navigator.  
Sök efter det önskade området och dra det till den cell i den aktuella tabellen där referensen skall infogas.  
Den här metoden kan du också använda om du vill infoga ett område från en annan tabell från samma dokument i den aktuella tabellen, d.v.s. i 3D-tabeller.  
Referenser till andra tabeller  
Du kan göra en referens till en cell i en annan tabell synlig i en tabellcell.  
Öppna ett nytt tomt tabelldokument.  
Mata in följande formel i t.ex. cell A1 i Tabell1 och avsluta inmatningen genom att trycka på returtangenten:  
=Tabell2.A1  
Om du nu klickar på tabellfliken med beteckningen Tabell2 vid undre fönsterkanten kommer du till Tabell2 i det aktuella dokumentet.  
Placera där markören i cell A1 och mata in en text eller ett tal.  
Om du växlar tillbaka till Tabell1, ser du där samma innehåll i cell A1.  
När innehållet i Tabell2.A1 ändras, ändras även innehållet i Tabell1.A1.  
En referens kan på motsvarande sätt också göras till en cell i ett annat dokument.  
Öppna ett annat dokument som redan är sparat som fil (detta fungerar inte med dokument som inte har sparats än).  
Om exemplen finns med i din installation kan du t.ex. öppna dokumentet Bio1 från tabellexemplen via kommandot Arkiv - Öppna.  
Placera markören i en tom cell och mata in ett likhetstecken som tecken på att du vill börja mata in en formel.  
Klicka där i cell C3.  
Växla tillbaka till det nya tabelldokumentet.  
På formellisten ser du nu hur %PRODUCTNAME Calc har kompletterat referensen i formeln åt dig.  
Där står till exempel nu:  
=' file: / //C_BAR_ / {installpath} / share / samples / swedish / spreadsheets / Bio1.sdc '#$Biobesök.C3  
Bekräfta formeln genom att klicka på den gröna bocken.  
Referensen till en cell i ett annat dokument innehåller alltså namnet på det andra dokumentet med enkla 'citattecken', sedan #-tecknet, sedan namnet på tabellen i det andra dokumentet följt av en punkt och namnet på cellen C3.  
Namnet på tabellen fick automatiskt ett ledande dollartecken, eftersom tabellen adresseras absolut.  
Om du undersöker namnet på det andra dokumentet i den här formeln ser du att det är skrivet som en URL.  
Om du nu tror att du kan ange en webbadress (URL) från Internet också, har du rätt.  
Om du t.ex. hittar en Internetsida med aktuella börskurser i tabellceller, kan du ladda den här sidan i %PRODUCTNAME Calc.  
Gör så här:  
Placera markören i den cell där du vill infoga externa data i ett %PRODUCTNAME Calc-dokument.  
Välj Infoga - Externa data.  
Dialogrutan Externa data visas.  
Mata in URL för ett dokument eller en webbsida i dialogrutan.  
Använd följande fullständiga URL-skrivsätt: (fiktivt exempel) http: / /www.min-bank.com / tabell.html.  
Du kan också mata in ett filnamn från det lokala filsystemet eller från ett nätverks filsystem på det här sättet, som i en Öppna-fil-dialogruta.  
%PRODUCTNAME laddar den angivna webbsidan eller filen "i bakgrunden", d.v.s. utan att visa den.  
I den stora listrutan i dialogrutan Externa data står namnen på alla tabeller eller områden som du nu kan välja ifrån.  
Välj ut en eller flera tabeller eller områden, aktivera den automatiska uppdateringen var n sekund om du vill och klicka på OK.  
Innehållet infogas som länk i %PRODUCTNAME Calc-dokumentet.  
Spara ditt tabelldokument.  
När du öppnar det igen senare kommer %PRODUCTNAME Calc att uppdatera innehållet i de länkade cellerna efter en bekräftelsefråga.  
Under Verktyg - Alternativ - Tabelldokument - Allmänt kan du välja att länkar i tabelldokumentet alltid, på begäran eller aldrig skall uppdateras automatiskt när du öppnar det.  
Uppdatering kan utlösas manuellt i dialogrutan Redigera - Länkar.  
Referera till en cell i ett annat dokument  
Du kan också referera till en cell i ett annat tabelldokument:  
Öppna ett tabelldokument där det redan finns ett innehåll eller mata in några tal och lite text i ett tabelldokument och spara det på hårddisken.  
Vi utgår i detta exempel från dokumentet 'C:\test\test.sxc' som innehåller en tabell med namnet Tabell1.  
Öppna ett nytt tomt tabelldokument  
Placera t.ex. markören i cell A1 och ange följande formel: =' C:\test\test.sxc '#Tabell1.A1  
Du kan även ange namnet på filen med URL-skrivsättet: =' file: / //C_BAR_ / test / test.sxc '#Tabell1.A1.  
Som du säkert förstår kan man referera till en fil på Internet på samma sätt, t.ex. 'http: / /www.sun.se / test / test.sxc'#Tabell1.A1 (fiktivt exempel).  
Om du nu utvidgar markeringen genom att dra i den lilla utvidgningsrutan i det nedre högra hörnet på den aktuella cellen, infogar %PRODUCTNAME de anpassade referenserna i de angränsande cellerna.  
Tabellnamnet används som absolut referens genom ett framförställt $-tecken.  
Tilldela format med formel  
Tillsammans med funktionen AKTUELL kan du ge cellen en viss färg beroende på vilket värde den innehåller.  
Annars får den cellformatmallen "Green".  
Om du vill utvidga samtliga celler i ett markerat område med en formeldel kan du använda dialogrutan Sök och ersätt.  
Markera alla celler som du vill utvidga.  
Välj kommandot Redigera - Sök och ersätt.  
Skriv följande i fältet Sök efter. .* (punkt asterisk)  
(.* är ett reguljärt uttryck som betecknar hela innehållet i den aktuella cellen.)  
Skriv följande i fältet Ersätt med: =&+FORMATMALL( OM(AKTUELL()>3 ;"Red" ;"Green"))  
(Tecknet & betecknar det aktuella innehållet i fältet Sök efter.  
I början på raden står likhetstecknet, eftersom vi vill infoga en formel.  
Vi utgår ifrån att de båda cellformatmallarna "Red" och "Green "redan finns.)  
Markera fälten Reguljärt uttryck och Bara markering.  
Klicka på Sök alla.  
Nu skall samtliga celler som fanns med i markeringen och som har ett innehåll vara framhävda.  
Klicka på Ersätt alla.  
Använda villkorlig formatering  
Med menykommandot Format - Villkorlig formatering kan du i en dialogruta definiera upp till tre villkor per cell som måste vara uppfyllda för att de markerade cellerna skall få ett visst format.  
På det här sättet kan du t.ex. i en cell med summor framhäva de summor som ligger över genomsnittet för samtliga summor.  
Om summorna ändras så ändras formateringen på motsvarande sätt utan att du behöver tilldela andra formatmallar manuellt.  
Markera de celler som skall få en villkorlig formatmall.  
Välj kommandot Format - Villkorlig formatering.  
Mata in villkoret / villkoren i den dialogruta som visas.  
Dialogrutan beskrivs utförligt i %PRODUCTNAME -hjälpen och nedan följer ett exempel på villkorlig formatering.  
Exempel på villkorlig formatering; skapa talvärden  
I en tabell med omsättningar kan du t.ex. lägga en grön bakgrund för alla värden som ligger över genomsnittet och en röd bakgrund för alla värden som ligger under.  
Detta kan du åstadkomma med den villkorliga formateringen.  
Fyll i en tabell med olika tal.  
Du kan skapa tabeller med slumptal:  
Du får då ett slumptal mellan 0 och 1.  
Om du vill ha heltal mellan 0 och 50 skriver du formeln =HELTAL( SLUMP()*50).  
Dra formeln till det önskade antalet celler i horisontell riktning.  
Muspekaren blir då ett hårkors.  
Håll ner musknappen och dra åt höger tills du har täckt önskat antal celler.  
Dra på samma sätt som är beskrivet ovan hörnet på cellen längst till höger nedåt, så att fler rader med slumptal skapas.  
Exempel på villkorlig formatering: definiera cellformatmallar  
I det här exemplet skapar du nu två cellformatmallar för dina tal: en mall för alla värden som visar omsättningar över genomsnittet och en för omsättningar som ligger under genomsnittet.  
Stylist bör nu vara synlig.  
Öppna snabbmenyn och välj Formatera celler.  
Klicka på fliken Bakgrund i dialogrutan Cellattribut och välj t.ex. ljusgrön som bakgrundsfärg.  
Klicka på OK.  
Klicka på ikonen Ny formatmall från markering i Stylist.  
Ge den nya mallen ett namn i dialogrutan, t.ex. "Över".  
För att definiera en andra mall klickar du återigen på en tom cell och gör som beskrivs ovan.  
Formatera cellen med bakgrundsfärgen ljusröd och kalla mallen för "Under".  
Exempel på villkorlig formatering: beräkna medelvärde  
I det här exemplet beräknas medelvärdet av slumptalen.  
Resultatet placeras i en cell:  
Placera cellmarkören i en tom cell, t.ex. J14, och starta funktionsautopiloten.  
Välj funktionen MEDEL.  
Markera samtliga slumptal med musen.  
Om funktionsautopiloten döljer området, kan du tillfälligt förminska dialogrutan med Förstora / Förminska.  
Stäng funktionsautopiloten med OK.  
Exempel på villkorlig formatering: använda cellformatmallar  
Nu behöver du bara använda den villkorliga formateringen på din tabell.  
Markera alla celler med slumptalen i tabellen.  
Välj kommandot Format - Villkorlig formatering....  
Dialogrutan Villkorlig formatering visas.  
Välj nu följande villkor:  
Om cellvärdet är mindre än J14, formatera då med "Under" och om cellvärdet är lika med eller större än J14, formatera då med "Över ".  
Exempel på villkorlig formatering: kopiera cellformatmallar  
Du vill använda den villkorliga formateringen på fler celler i efterhand:  
Klicka på en av cellerna som har villkorlig formatering.  
Kopiera cellen till urklippet, t.ex. med Kommando Ctrl +C.  
Markera cellerna som ska ha samma formatering.  
Välj kommandot Redigera - Klistra in innehåll.  
Dialogrutan Klistra in innehåll.  
Markera bara fältet Format i området Urval, avmarkera de andra.  
Klicka på OK.  
Format - Villkorlig formatering  
Framhäva negativt tal  
Du kan också definiera ett eget talformat där negativa tal framhävs med andra färger.  
Markera cellerna och välj kommandot Format - Cell.  
Klicka på fliken Tal, välj ett talformat och markera rutan Negativa värden i rött.  
Klicka på OK.  
Cellerna får ett talformat vars formatkod är definierad i två delar.  
Efter semikolonet står formatet för negativa tal.  
Koden [RED] kan du ändra i textfältet Formatbeskrivning.  
Mata t.ex. in YELLOW istället för RED.  
När du infogat den nya koden i listan genom att klicka på ikonen Lägg till har du matat in en giltig färgkod.  
Använda cellformatmallar  
Öppna ett nytt tomt tabelldokument.  
Placera markören i cell A1 och skriv in en text.  
Placera markören i cell A2 och skriv in ett tal.  
Formatera talet som resultat genom att tilldela det cellformatmallen "Resultat".  
Placera markören i cellen, visa Stylist (F11) och dubbelklicka sedan på posten "Resultat ".  
Formatera texten som överskrift med till exempel fet stil, 20 punkters storlek och blå text på gul bakgrund.  
Placera markören i A1, mata in de önskade attributen med ikonerna och listrutorna på textobjektlisten.  
Du kan också markera hela texten i cellen och sedan öppna snabbmenyn till den markerade texten och välja kommandot Tecken.  
Det här nya formatet skall nu definieras som ny formatmall.  
Klicka på symbolen Ny formatmall från markeringen i Stylist.  
En dialogruta visas där du kan skriva ett namn på den nya formatmallen.  
Du kan t.ex. kalla den nya cellformatmallen för "Rubrikformat".  
Klicka på OK.  
Den nya cellformatmallen visas i Stylist.  
Om du vill tilldela celler det nya rubrikformatet, markerar du dem och dubbelklickar på cellformatmallens namn i Stylist.  
Upphäva cellskydd  
Gå till tabellen, vars skydd du vill upphäva.  
Du väljer Verktyg - Skydda dokument, klickar sedan antingen på Tabell eller Dokument för att upphäva markeringen.  
Om du har lämnat ett lösenord måste du nu ange det i en dialogruta och bekräfta dialogrutan med OK.  
Cellerna kan nu redigeras, formlerna kan göras synliga och alla celler skrivas ut igen, tills du aktiverar skyddet för tabellen eller dokumentet på nytt.  
Konsolidering av data  
Vid konsolidering sammanfogas cellinnehållet från flera tabeller i det aktuella dokumentet på ett ställe.  
Du väljer en beräkningsregel så att t.ex. summan, standardavvikelsen eller variansen för data visas i konsolideringsområdet.  
1.  
Växla till dokumentet med områdena som ska konsolideras.  
2.  
Välj dialogrutan Data - Konsolidera.  
Dialogrutan Konsolidera visas.  
3.  
I listrutan Källdataområde väljer du ett område som du vill utgå ifrån och sammanfoga med andra områden.  
4.  
Om området inte har något namn, klickar du i inmatningsfältet till höger om listrutan Källdataområde.  
Då ser du en blinkande textmarkör där.  
Skriv nu referensen till det första källdataområdet med tangentbordet, eller markera det med musen i tabellen.  
5.  
Klicka på Lägg till för att lägga till det markerade området i fältet Konsolideringsområden.  
Området visas där.  
6.  
Välj nu ut ytterligare områden med en av de beskrivna metoderna, och klicka på Lägg till efter varje område.  
7.  
Bestäm var resultatet ska matas ut genom att markera målområdet i listrutan Resultat vid.  
8.  
Använd tangentbordet till att skriva in områdesadressen till målområdet eller adressen till den vänstra övre cellen i målområdet.  
Alternativt kan du också markera målområdet med musen eller sätta cellmarkören i målområdets vänstra övre cell.  
9.  
Välj en beräkningsregel, enligt vilken konsolideringsområdenas värden ska sammankopplas med varandra.  
Summafunktionen är förinställd för enkel addition av alla värden som hör samman.  
10.  
Klicka på OK om du vill konsolidera områdena.  
Om du inte vill skapa en ny tabell som är oberoende av utgångsområdena utan en tabell där länkarna till källområdena finns kvar, eller om du vill sammanfoga områden där ordningsföljden för rader eller kolumner är olika, klickar du på Fler.  
Dialogrutan Konsolidera utvidgas.  
Nu placeras inte resultaten av beräkningen som värden i konsolideringens målområde, utan formlerna som har lett till dessa resultat.  
På det här sättet kommer en ändring i efterhand i ett av källområdena också att ändra det tillhörande målområdet.  
Dessa rader delas in automatiskt och döljs, och bara slutresultatet visas på en rad enligt den valda beräkningsregeln.  
Nu sammanfogas cellerna i källområdena inte 1:1 enligt cellens position i området, utan enligt samma radetikett eller samma text i kolumnhuvudena.  
De här texterna måste markeras med musen när källområdena markeras.  
Texterna måste vara identiska, så att raderna eller kolumnerna tilldelas korrekt.  
Om skrivsättet i en rad eller kolumn avviker från de andra, bifogas den i slutet av målområdet som ny rad eller kolumn.  
Konsoliderings - och målområdenas data sparas.  
När du öppnar ett dokument där en konsolidering har definierats, står dessa data till förfogande igen.  
Data - Konsolidera  
Formler och värden som csv-fil  
Csv-filer är rena textfiler där cellinnehåll från en tabell finns.  
Som fältavgränsare mellan cellerna används t.ex. komma eller semikolon.  
Texter sätts automatiskt inom citationstecken, tal skrivs direkt.  
Export av formler och värden som csv-fil  
Växla till tabellen som ska skrivas som csv-fil.  
Om du vill exportera formlerna som formler, t.ex. i form av =SUMMA( A1:B5), gör du så här:  
Välj Verktyg - Alternativ - Tabelldokument - Vy.  
I området Visa markerar du rutan Formler.  
Klicka på OK.  
Om du vill exportera de beräknade resultaten i stället för formlerna, får inte rutan Formler vara markerad.  
Välj Arkiv - Spara som.  
Dialogrutan Spara som öppnas.  
I fältet Filtyp väljer du formatet "Text CSV".  
Ange ett namn och klicka på Spara.  
I dialogrutan Textexport som öppnas väljer du teckenuppsättningen samt fält - och textavgränsare för de data som ska exporteras och bekräftar med OK.  
OBS:  
Om talen innehåller komman som decimaltecken eller tusentalsavgränsare, får du inte välja komma som fältavgränsare!  
Om det finns dubbla citattecken i texterna måste du välja enkelt citattecken (apostrof) som textavgränsare och tvärtom.  
Avmarkera eventuellt rutan Formler igen när du har sparat så att du ser de beräknade resultaten i tabellen igen.  
Import av en csv-fil  
Välj Arkiv - Öppna.  
Dialogrutan Öppna visas.  
I fältet Filtyp väljer du formatet "Text CSV".  
Välj filen och klicka på Öppna.  
Om filen har .csv som filnamnstillägg, identifieras filtypen automatiskt.  
Dialogrutan Textimport öppnas.  
Klicka på OK.  
Om csv-filen innehåller formler som formler, avmarkerar du rutan Formler (i Verktyg - Alternativ - Tabelldokument - Vy) så att du ser de beräknade resultaten i tabellen.  
Verktyg - Alternativ - Tabelldokument - Vy  
Textexport  
Textimport  
Celler i valutaformat  
Om du klickar på ikonen Talformat: valuta på objektlisten för att formatera ett tal, får cellen det standardvalutaformat som är inställt under Verktyg - Alternativ - Språkinställningar - Språk i %PRODUCTNAME.  
Detta kan leda till missförstånd vid internationellt utbyte av %PRODUCTNAME Calc-dokument.  
Tänk dig att ditt %PRODUCTNAME Calc-dokument laddas av en annan användare som använder ett annat standardvalutaformat.  
I %PRODUCTNAME Calc kan du definiera att ett tal som du t.ex. har formaterat som "1 234,50 €" anges som euro även i ett annat land och inte som t.ex. dollar.  
Du kan påverka valutaformatet i dialogrutan Cellattribut (meny Format - Cell - flik Tal) med två landsinställningar.  
I listrutan Språk väljer du grundinställningen för valutatecken, decimaltecken och tusentalsavgränsare.  
I listrutan Format väljer du eventuella avvikelser i valutatecknet från formatet som definieras genom språket.  
Om språket till exempel är inställt till "Standard" och du använder en tysk språkvariant, är valutaformatet "1.234,00 €".  
För att gruppera siffrorna i tusental används punkt och framför decimalerna ett komma.  
Om du väljer "$Engelska (US)" som valutaformat i listrutan Format får du följande format: "$ 1.234,00 ".  
Som du ser är decimaltecknen desamma.  
Bara valutatecknet har ändrats och placerats om, men formatet som ligger till grund för talets skrivsätt är så som det har definierats genom språkvarianten.  
Om du ställer om språket för cellerna till "Engelska (US)" från början, används även den engelska språkvarianten för avgränsarna och standardformat för valuta är nu "$ 1,234.00 ".  
Även här kan du ändra formatet, t.ex. till "1,234.00 €".  
Det här skrivsättet för tal är mer bekant för en användare av ett amerikanskt system.  
Format - Cell - Tal  
Definiera databasområde  
Om du till exempel vill administrera dina hushållskostnader elektroniskt, kan du mata in dataposterna i ett nytt %PRODUCTNAME Calc-tabelldokument och definiera området som databasområde.  
Skapa dataposter i tabelldokument  
Öppna ett nytt, tomt tabelldokument.  
Skriv rubriken för kolumnerna på den första raden, t.ex. "Datum" i cell A1, "Användning "i B1, "Belopp" i C1 och mata in lite data.  
Om du vill formatera din tabell som på bilden gör du så här:  
1.  
Markera rad 1 genom att klicka på radhuvudet.  
Klicka på ikonen Fet.  
2.  
Markera hela kolumn A genom att klicka på kolumnhuvudet.  
Öppna snabbmenyn och välj Formatera celler.  
Välj ett datumformat för kolumn A som det visas på bilden.  
3.  
Markera hela kolumn C genom att klicka på kolumnhuvudet och tilldela den ett valutaformat.  
Det räcker att klicka på ikonen Talformat: valuta på objektlisten.  
Definiera databasområde  
Definiera det markerade området som %PRODUCTNAME Calc-databasområde genom att välja Data - Definiera område.  
I dialogrutan Definiera databasområde är det markerade området redan registrerat.  
Markera i varje fall rutan Innehåller kolumnhuvuden så att den första raden kommer med.  
Den här rutan visas om du klickar på Fler.  
Mata in ett namn på området och stäng dialogrutan med OK.  
Nu har du definierat det markerade området som databasområde, vilket bland annat innebär att du lätt kan sortera raderna (= dataposterna).  
Sorteringar, filtreringar o.s.v. som du har definierat för databasområdet uppdateras.  
Filtrera databasområde  
Om du bara vill filtrera fram vissa dataposter från längre datalistor för att fortsätta att redigera dem, så kan du använda filterfunktionerna i tabelldokument.  
Du kan välja mellan att antingen definiera kriterierna exakt i en dialogruta där även områdesdefinitioner är möjliga eller att skapa ett AutoFilter som sedan alltid hjälper dig när du vill filtrera efter bestämda värden eller texter.  
Tänk dig till att börja med att utgiftslistan har mer än 8000 dataposter.  
Då kan du inte längre överblicka den själv.  
Nu vill du bara se dataposterna som har tillkommit efter den 2 / 1/2000 och som dessutom har ett belopp på över 500 valutaenheter.  
Placera markören i databasområdet och välj Data - Filter - Standardfilter.  
Mata in följande: datum > 2 / 1/2000 OCH belopp > 500.  
Som du ser kan du lätt välja ut datafältens innehåll i kombinationsfälten, men du kan också mata in beloppet 500 direkt.  
När du klickar på OK ser du bara dataposterna som uppfyller alla kriterier.  
Återställ visningen igen med menykommandot Data-Filter-Ta bort filter.  
Om du bara vill visa dataposter som har ett bestämt innehåll är det lätt att använda AutoFilter:  
Placera markören i databasområdet.  
Klicka på ikonen Automatiskt filter på verktygslisten.  
Nu har kolumnhuvudena i databasområdet fått små kommandoknappar.  
Klicka på kommandoknappen bredvid Datum och välj till exempel 00-01-02.  
Du ser bara dataposterna med det här datumet.  
Genom att klicka på ikonen Automatiskt filter på verktygslisten återställer du visningen igen.  
Gruppera databasområde och beräkna delsummor  
Om du vill utöka exempeluppgifterna och använda dem som hushållsbudget vill du säkert också sammanfatta och skriva ut utgifterna i del - och slutresultat.  
Även detta är möjligt med några få steg.  
Placera markören i databasområdet.  
Välj Data - Delresultat.  
Du ser dialogrutan Delresultat.  
Mata in de önskade alternativen för beräkning av delsummor:  
Gruppera delresultat efter "Datum" (det innebär att en ny delsumma beräknas så snart ett nytt datum börjar) och beräkna dem för "Belopp "med beräkningsregeln "Summa" (alltså summera delresultatens belopp).  
Så snart du trycker på returtangenten eller klickar på OK ser du effekterna: tabellen grupperas efter delresultat.  
Den totala summan visas längst ner.  
Lägg märke till styrelementen till vänster om radhuvudena.  
Där kan du se igen vilka dataposter (= rader) som har sammanfattats.  
Om du klickar på ett minustecken visas bara den sammanfattande resultatraden.  
Men det är enklast att styra strukturen med de små siffrorna i övre kanten av grupperingsområdet.  
Om du klickar på den lilla 1:an, så ser du bara den totala summan; 2:an visar dessutom delsummorna och 3:an visar allt.  
Sortera databasområde  
Du har markerat ett cellområde och definierar det som databasområde med Data - Definiera område.  
Placera markören i databasområdet och öppna dialogrutan Data - Sortera.  
Där väljer du kolumnen som ska sorteras, t.ex. "Belopp", som sorteringskriterium och klickar på OK.  
Du kan ange upp till ytterligare två underordnade sorteringskriterier, till exempel först sortera utgifterna efter datum, vid samma datum efter post och vid samma datum och post efter belopp.  
Skapa datapilottabell  
Markera dataområdet för en tabell tillsammans med rad - och kolumnhuvudena.  
Välj Data - Datapilot - Starta.  
Dialogrutan Välj ut källa visas.  
Välj alternativet Aktuell markering och bekräfta med OK.  
I dialogrutan Datapilot visas tabellens kolumnhuvuden som kommandoknappar, som du fritt kan placera med hjälp av dra-och-släpp i layoutområdena "Kolumn", "Rad" och "Data ".  
Dra önskade fält till ett av de tre områdena.  
Fältet placeras där.  
Om kommandoknappen placeras i området Data får det en etikett som även visar formeln som används för att skapa data i dataområdet.  
Genom att dubbelklicka på ett av fälten i området Data öppnar du dialogrutan Datafält.  
Här kan du välja den funktion som används för visning av data i dataområdet.  
Du kan välja flera funktioner genom att hålla ner Ctrl-tangenten när du klickar med musen.  
Du kan när som helst ändra ordningsföljden på kommandoknapparna genom att flytta dem inom området med musen.  
Du lägger tillbaka en kommandoknapp genom att flytta den från området till de andra kommandoknapparna med musen.  
Om du dubbelklickar på en av kommandoknapparna i området Rad eller Kolumn, öppnas dialogrutan Datafält.  
Här kan du välja om och i vilken omfattning %PRODUCTNAME ska räkna ut och visa delresultat.  
Avsluta datapiloten med OK.  
I tabellen infogas nu - standardpositionen är under det markerade området - en kommandoknapp som heter Filter och två rader längre ned den beräknade datapilottabellen.  
Den är omgiven av en tjock linje.  
Radera datapilottabell  
Sedan väljer du Data - Datapilot - Radera.  
Redigera datapilottabell  
Klicka på en av kommandoknapparna i tabellen som datapiloten har skapat och håll ner musknappen.  
Vid muspekaren visas en särskild symbol.  
Dra kommandoknappen till en annan position på raden om du vill ändra kolumnernas ordningsföljd.  
Dra kommandoknappen från raden i tabellens vänstra kant till radhuvudenas område, om du vill göra en rad av en kolumn.  
Muspekaren ändrar sitt utseende från symbol för kolumnhuvud till symbol för radhuvud.  
Om du vill ta bort en kommandoknapp från tabellen drar du ut den från tabellen.  
Släpp musknappen när muspekaren har förvandlats till ett förbudstecken på tabellarket.  
Kommandoknappen är då raderad.  
Om du dubbelklickar på namnet på ett tabellelement visas respektive döljs de element som finns under det.  
Filtrera datapilottabell  
Även om datapilottabellen i regel skapas efter användarens önskemål, kan det förekomma att inte alla data som finns i tabellen är av intresse.  
I sådana fall använder man filter, som med hjälp av vissa villkor filtrerar bort motsvarande data från den befintliga tabellen.  
Du öppnar inmatningsmasken för filtervillkoren genom att klicka på kommandoknappen Filter i datapilottabellen på tabellarket.  
Du ser dialogrutan Filter.  
Den här dialogrutan innehåller olika kriterier för dataurval.  
Välja utdataområde för datapilottabell  
Klicka på kommandoknappen Fler i dialogrutan Datapilot.  
Dialogrutan utvidgas.  
I listrutan Utdata från kan du välja ett område försett med namn, där datapilottabellen ska skapas.  
Om utdataområdet inte har något namn, anger du adressen för områdets övre vänstra cell i fältet till höger om listrutan Utdata från.  
Du kan också klicka med musen på cellen för att mata in cellens adress här.  
Om du kryssar för rutan Ignorera tomma rader, tas inte hänsyn till tomma rader när datapilottabellen skapas.  
Om du kryssar för rutan Identifiera kategorier, identifieras och tilldelas kategorier med hjälp av överskrifterna när datapilottabellen skapas.  
Uppdatera datapilottabell  
Om data i grundtabellen ändras, måste %PRODUCTNAME genomföra beräkningen av tabellen på nytt för att uppdatera utvärderingen.  
Om du vill genomföra en ny beräkning i tabellen, håller du ner Ctrl-tangenten höger musknapp och klickar på ett av kommandoknappfälten och väljer Uppdatera eller Data - Datapilot - Uppdatera.  
Datapilot  
Datapiloten ger dig möjlighet att analysera och utvärdera redan inmatade data.  
Den gör det möjligt att skapa olika rapporter utifrån samma värden, beroende på vilken aspekt som står i förgrunden för analysen.  
Tänk dig t.ex. en dataanalystabell som innehåller ditt företags försäljningsdata, för vissa varugrupper, filialer och år.  
Med hjälp av datapiloten kan du alltid snabbt genomsöka tabellen efter aktuella, intressanta data.  
Vad behöver du datapiloten till?  
En tabell som är skapad med hjälp av datapiloten är en interaktiv tabell, vilket innebär att data kan ordnas, omordnas eller sammanfattas utifrån olika aspekter.  
Denna funktion är tillämplig t.ex. vid försäljningsstyrning.  
För det första kan det vara viktigt att studera omsättningssiffrorna inom en viss tidsram, för det andra kan det vara relevant att utvärdera försäljningssiffrorna efter regionala aspekter.  
Temaurval för en tabell  
Det bästa är att öppna ett av de exempeldokument som finns i mappen Exempel - Tabeller i %PRODUCTNAME.  
De här exempeltabellerna har skapats med de utbytbara användarformatmallarna.  
Du kan öppna Stylist och ställa in vyn på användarformatmallarna i den nedre listrutan.  
Nu ser du en lista över de användardefinierade cellformatmallar som finns i det aktuella dokumentet.  
Så snart du väljer ett annat tema i dialogrutan Temaurval byts några av egenskaperna i användarformatmallarna ut.  
Ändringarna visas omedelbart i tabellen, i den mån respektive användarformatmall har tilldelats tabellen.  
När du skapar ett eget tabelldokument, kan du förse det med utbytbara användarformatmallar.  
Användarformatmallarna finns nu till hands och syns i Stylist.  
Genom att dubbelklicka på en användarformatmalls namn i Stylist kan du använda formatmallen på de markerade cellerna.  
Temaurval  
Kalkera flera tabeller  
Du vill ange nya likadana kolumn - och radrubriker för alla tre tabellerna.  
Markera alla tre tabellerna genom att hålla ner skifttangenten och klicka på alla gråa registerflikar i nedre kanten av arbetsområdet.  
Sedan är alla tre registerflikar vita.  
De visas sedan i samma position även i de andra markerade tabellerna.  
Räkna om eurobelopp med formel  
Om du vill räkna om 500 kr till euro kan du skriva följande formel i en cell:  
=OMRÄKNA( 500 ;"SEK" ;"EUR")  
Som resultat får du antalet euro för 500 kronor.  
Beloppet som ska omräknas står alltså alltid först i parentesen.  
Det kan anges direkt, som här, eller som referens.  
Om t.ex. beloppet står i cell D2 kan du ange D2 som första del av funktionen i formeln.  
De andra delarna i funktionen är beloppets enhet och enheten som beloppet ska omräknas till.  
Alla tre delarna i funktionen avgränsas med semikolon.  
Med formeln =OMRÄKNA( 50 ;"EUR" ;"SEK") får du veta hur många kronor 50 euro är värda.  
Om du har ett antal SEK-belopp under varandra i kolumn D från D2 till D20 och vill ha samma belopp i euro i kolumn E från E2 till E20, gör du så här:  
Klicka i cell E2.  
Mata in följande: =OMRÄKNA (  
Klicka i cell D2.  
Nu är D2 definierad som första del av funktionen.  
Markören står fortfarande på D2 i formeln.  
Mata in följande text:; "SEK" ;"EUR "  
(skriv texten med båda semikolon och citationstecknen) och tryck på returtangenten.  
Därmed är hela formeln avslutad; den lyder =OMRÄKNA(D2 ;"SEK" ;"EUR").  
I cellen E2 står nu resultatet av beräkningen.  
Klicka i cell E2, sedan i den lilla kvadraten längst ner till höger i cell E2 och håll ner musknappen och dra neråt till cell E20.  
Släpp musknappen där.  
Nu har du kopierat formeln från E2 till E20.  
Referenserna har automatiskt anpassas så att de alltid hänvisar till den angränsande cellen till vänster.  
AutoPilot Eurokonverterare  
Använda filter  
Med hjälp av filter och specialfilter kan du uppnå att bara vissa rader = dataposter i ett dataområde är synliga.  
I tabelldokumenten i %PRODUCTNAME finns det flera möjligheter att använda filter.  
Du kan använda AutoFilter -funktionen för att bara visa de dataposter som har samma post i ett datafält.  
Med hjälp av filterdialogrutan kan du dessutom definiera gränser för värdena, så att bara de dataposter visas vars värden ligger inom de definierade gränserna.  
Du kan kombinera upp till tre villkor av detta slag med logiskt OCH eller logiskt ELLER.  
Detta är standardfiltret.  
Specialfiltret slutligen går utöver denna begränsning på tre villkor och medger sammanlagt upp till åtta filtervillkor.  
Med specialfilter skriver du in villkoren direkt i tabellen.  
Om du markerar några rader med filter och sedan vill radera dem, måste du först hålla ner Ctrl-tangenten och klicka på alla rader som är synliga efter filtreringen innan de raderas.  
Då kan du vara säker på att bara de raderna är markerade och att bara de raderas.  
Utforma tabelldokument översiktligt  
I %PRODUCTNAME finns det ett flertal möjligheter att utforma tabeller snabbt utan mycket arbete.  
Som exempel visar vi här tre olika versioner av samma tabell som bara skiljer sig åt i formateringen:  
Här ser du en exempeltabell utan någon formatering, vilket motsvarar standardutseendet.  
Om samma tabell bara formateras med ett av AutoFormaten får man utan vidare efterbearbetning en snygg bild.  
Här har exempeltabellen formaterats med några cellattribut i dialogrutan Format - Cell.  
Dessutom har visningen av gitterlinjer och tabellhuvuden tagits bort via Verktyg - Alternativ - Tabelldokument - Vy och en grafikfil har laddats som bakgrundsbild via Format - Sida - Bakgrund.  
En bild som du laddar via Format - Sida - Bakgrund är bara synlig på en utskrift och via menykommandot Arkiv - Förhandsgranskning.  
Om du vill ha en bakgrundsbild även på bildskärmen, infogar du ett grafikobjekt via Infoga - Grafik - Från fil och placerar sedan grafikobjektet bakom cellerna via snabbmenykommandot Placering - I bakgrunden.  
Använd Navigator om du vill markera det här grafikobjektet i bakgrunden igen senare.  
Så här formaterar du text i ett tabelldokument  
Markera texten som du vill formatera.  
Välj textattributen på tabellobjektlisten eller välj Format - Cell.  
Du ser då dialogrutan Cellattribut där du kan välja textattribut, framför allt under fliken Teckensnitt.  
Så här formaterar du talvisningen i ett tabelldokument  
Markera cellerna där du vill ändra talvisning.  
Om du vill formatera talen i standard-valutaformat eller som procenttal hittar du motsvarande ikoner på tabellobjektlisten.  
För andra format väljer du Format - Cell.  
Under fliken Tal kan du välja ut formaten och definiera egna format.  
Så här formaterar du kanter och bakgrund för celler och sidor  
Som regel gäller att du kan tilldela varje grupp av celler ett format genom att först markera cellerna (om du håller ner Kommandotangenten Ctrl-tangenten kan du göra multimarkeringar) och sedan öppna dialogrutan Cellattribut via Format - Cell.  
Välj sedan till exempel inramning och bakgrund.  
Om du vill formatera hela utskriftssidan väljer du Format - Sida.  
Du kan sedan till exempel mata in sidhuvud och sidfot som visas på varje sida vid utskrift.  
Formatera tal  
Mata in ett tal i tabellen, till exempel 1234,5678.  
Du ser därför 1234,57 när du bekräftar din inmatning.  
Men internt behåller talet sina fyra decimaler efter decimaltecknet och avrundas bara när det visas i dokumentet.  
Placera markören på talet och öppna nu dialogrutan Cellattribut genom att välja Format - Cell.  
Nu ser du ett urval av talformat.  
Nere till höger i dialogrutan ser du en förhandsvisning av hur ditt aktuella tal skulle se ut om du väljer ett visst format.  
I dialogrutan kan du förutom talformaten också bestämma andra attribut som skall gälla för de markerade cellerna eller det markerade cellinnehållet.  
Under fliken Teckensnitt kan du t.ex. definiera teckensnitt, -storlek och -färg.  
Om du bara vill ändra antalet visade decimaler är det enklast att använda ikonen Talformat: lägg till decimal respektive Talformat: radera decimal på objektlisten.  
Kopiera formel  
Det finns flera sätt att kopiera en formel, gör t.ex. så här:  
Markera cellen som innehåller formeln.  
Välj Redigera - Kopiera.  
Du kan också använda tangentkombinationen Kommando Ctrl +C för kopiering.  
Markera cellen som formeln skall kopieras till.  
Välj Redigera - Klistra in eller använd tangentkombinationen Kommando Ctrl +V.  
Formeln anpassas korrekt i den nya cellen.  
Det finns ett mycket enkelt och snabbt sätt att kopiera till angränsande cellområden om du vill kopiera en formel till flera celler:  
Markera cellen som innehåller formeln.  
Klicka nere till höger i den framhävda ramen som omger cellen och håll ner musknappen.  
Muspekaren blir till ett hårkors.  
Dra neråt eller till höger med nertryckt musknapp över cellerna som du vill kopiera formeln till.  
Släpp musknappen.  
Formeln kopieras till cellerna och anpassas automatiskt korrekt.  
Om värden och texter inte skall anpassas automatiskt, håller du ner Kommandotangenten Ctrl-tangenten samtidigt som du drar med musen.  
Formler anpassas alltid.  
Mata in formel på formellisten  
Klicka på cellen där du vill mata in formeln.  
Klicka på ikonen Funktion på formellisten.  
Du ser nu ett likhetstecken på inmatningsraden och kan börja att mata in formeln.  
Avsluta inmatningen genom att trycka på Retur eller klicka på ikonen Överta.  
Om du vill avbryta inmatningen och ignorera innehållet på inmatningsraden trycker du på Esc eller klickar på ikonen Ignorera.  
Du kan naturligtvis skriva in värden och formler direkt i cellerna, även om inmatningsmarkören inte syns där.  
Formler måste alltid börja med ett likhetstecken.  
När du redigerar en formel med referenser, framhävs referenserna i formeln och de tillhörande cellerna i tabellen i samma färg.  
Då anpassas även referensen i formeln på inmatningsraden.  
Du kan stänga av Visa referenser i färg under Verktyg - Alternativ - Tabelldokument - Vy.  
Om du vill se en beräkning av de enskilda delarna i en sammansatt formel, så markerar du de enskilda delarna och trycker på F9.  
I formeln =SUMMA( A1:B12)*SUMMA(C1:D12) kan du t.ex. markera delen SUMMA(C1:D12) och trycka på F9.  
Då visas delresultatet i tipshjälpen.  
Om det blir fel i formeln du skapar visas en felkod i den aktiva cellen.  
Formellist  
Räkna med formler  
Alla formler börjar med ett likhetstecken.  
Även andra element är möjliga, som till exempel formatangivelser som bestämmer hur talen skall formateras.  
Formler kan naturligtvis också innehålla räkneoperatorer, logiska operatorer eller funktioner.  
Tänk på att även de fyra räknesätten kan användas med sina formeltecken +, -, * och / i formler, enligt regeln "punkträkning före streckräkning".  
I stället för =SUMMA( A1:B1) kan du skriva: =A1+B1.  
Även parenteser är möjliga.  
Formeln =1+2*3 returnerar något annat än =( 1+2 )*3.  
Här följer några exempel på %PRODUCTNAME Calc-formler:  
=A1+10  
Visar innehållet i A1 plus 10.  
=A1*16%  
Visar 16 procent av innehållet i A1.  
=A1 * A2  
Visar resultatet av multiplikation i A1 och A2.  
=AVRUNDA( A1;1)  
Avrundar innehållet i A1 till en decimal.  
=EFFRÄNTA( 5%;12)  
Beräknar effektiv ränta på 5% årligen och 12 betalningar.  
=B8-SUMMA( B10:B14)  
Beräknar summan av B10 till B14 och subtraherar värdet från B8.  
=SUMMA( B8;SUMMA(B10:B14))  
Beräknar summan av B10 till B14 och adderar värdet till B8.  
Du kan även skjuta in funktioner i formlerna som visas i exemplet.  
I stället för =AVRUNDA( A1;1) kan du alltså till exempel även beräkna formeln =AVRUNDA(SIN(A1);2).  
Funktionsautopiloten hjälper dig vid inskjutna funktioner.  
Lista med funktioner  
Funktionsautopilot  
Visa formler eller värden  
Om du vill visa formler i celler, t.ex. i form av =SUMMA( A1:B5), gör du så här:  
Välj Verktyg - Alternativ - Tabelldokument - Vy.  
I området Visa markerar du rutan Formler.  
Klicka på OK.  
Om du vill se de beräknade resultaten i stället för formlerna får rutan Formler inte vara markerad.  
Verktyg - Alternativ - Tabelldokument - Vy  
Mata in bråk  
Du kan även ange ett bråk i en cell och räkna med det:  
Mata in "0 1 / 5" i en cell (utan citationstecknen) och tryck på returtangenten.  
På inmatningsraden ser du värdet 0,2 som används för beräkningen.  
Om du skriver "0 1 / 2" ersätter AutoKorrigeringen de tre tecknen 1, / och 2 med ett enskilt tecken.  
Liknande gäller för 1 / 4 och 3 / 4.  
Den här ersättningen definieras under meny Verktyg - AutoKorrigering, fliken Ersättning.  
Om du vill kunna se flersiffriga bråk som "1 / 10", måste du ställa om cellformatet till visningen flersiffriga bråk (snabbmeny till cellen, kommando Formatera celler).  
Du kan sedan ange bråken 12 / 31 eller 12 / 32 - men bråken kortas automatiskt av så att du skulle se 3 / 8 i det sista exemplet.  
Använda målvärdessökning  
Med hjälp av målvärdessökning fastställer du ett värde, vilket som del av en formel leder till ett resultat som du fördefinierar av formeln.  
Du definierar alltså formeln med flera fasta värden och ett variabelt värde och resultatet av formeln.  
Det är lättast att förklara målvärdessökning med hjälp av ett exempel.  
För att beräkna den årliga räntan skapar du en tabell, som av värdena för kapital (K), antal år (i) och räntesatsen (p) ger resultatet - räntebelopp per år (R).  
Formeln lyder:  
R = K * i * p / 100  
Ränteintäkt = kapital * år * räntesats / 100.  
Sedan använder du variabelnamnen i följande exempel, d.v.s. namnet kapital istället för K o.s.v.  
I exemplet beräknas först att ränteinkomsten uppgår till 11 250 €per år med ett placerat kapital på 150 000 €och en räntesats på 7,5%. (Cellerna har formaterats i efterhand, A5 och E5 med valutaformat, C5 med procentformat.  
Sedan har cellbredderna anpassats.)  
Det är bäst att ge cellerna namn så att de kan användas med namn i formeln.  
Namnge celler  
Markera cell A5 i vårt exempel, sedan väljer du Infoga - Namn - Definiera.  
Dialogrutan Definiera namn visas.  
Skriv namnet K i textfältet.  
Längst ner i dialogrutan ser du referensen $Tabell1.$A$5 som du kan kontrollera.  
Klicka på Lägg till.  
Skriv in nästa namn i textfältet, sätt cellmarkören i cell B5 och klicka åter på Lägg till.  
Skriv in p i textfältet, sätt cellmarkören i cell C5 och klicka på Lägg till igen.  
Stäng dialogrutan med OK.  
Du kan nu också skriva formeln i E5 som = K * i * p istället för som =A5*B5*C5.  
Starta målvärdessökning  
Men vi undrar hur mycket kapitalinsatsen måste ändras för att vi ska uppnå en viss årsintäkt.  
Vi ska räkna ut hur mycket kapital som är nödvändigt för att ränteinkomsten ska uppgå till 15 000 €.  
Sätt markören i fältet E5 i tabellen.  
Välj Verktyg - Målvärdessökning.  
Dialogrutan Målvärdessökning visas.  
I fältet Formelcell är redan rätt cell angiven.  
Sätt markören i fältet Variabel cell i dialogrutan.  
A5, och klicka på den.  
Ange det önskade målvärdet, resultatet av formeln, i textfältet Målvärde i dialogrutan, i detta exempel 15000.  
Klicka på OK.  
Du får nu se en dialogruta som talar om att målvärdessökningen lyckats.  
Resultatet anges och om du vill kan du överta det.  
Klicka på Ja.  
Resultatet förs in i A5.  
Målvärdessökning  
Spara och öppna tabell som HTML  
Spara tabell som HTML  
%PRODUCTNAME Calc sparar alla tabeller i ett Calc-dokument tillsammans som HTML-dokument.  
I början av HTML-dokumentet infogas automatiskt en överskrift och en lista med hyperlänkar som leder till de olika tabellerna i dokumentet.  
Tal skrivs som visat.  
Dessutom skrivs det exakta interna värdet i HTML-taggen <SDVAL> så att du kan räkna med de exakta värdena när du har öppnat HTML-dokumentet med %PRODUCTNAME.  
Om du vill spara det aktuella Calc-dokumentet som HTML väljer du Arkiv - Spara som.  
Välj Filtyp "Webbsida".  
Ange ett Filnamn och klicka på Spara.  
Öppna tabell som HTML  
HTML-dokument öppnas alltid skrivskyddat.  
Om du vill redigera ett öppet HTML-dokument klickar du på ikonen Redigera fil på funktionslisten.  
%PRODUCTNAME har olika filter som du kan använda när du öppnar HTML-filer.  
Du väljer filter i dialogrutan Arkiv - Öppna i fältet Filtyp (lägg märke till området eftersom namnet "Webbsida "alltid är detsamma):  
Öppna i %PRODUCTNAME Writer / Web-filtret "Webbsida" eller med standardinställningen, d.v.s. utan att välja ett filter.  
Du har tillgång till alla möjligheter i %PRODUCTNAME Writer / Web, t.ex. kommandot Visa HTML-källtext.  
Öppna i %PRODUCTNAME Writer-filtret "Webbsida".  
Du har tillgång till alla möjligheter i %PRODUCTNAME.  
Men alla redigeringsmöjligheter som %PRODUCTNAME Writer har för dokument kan inte sparas i HTML-format.  
Öppna i %PRODUCTNAME Calc-filtret "Webbsida".  
Du har tillgång till alla möjligheter i %PRODUCTNAME Calc.  
Men alla redigeringsmöjligheter som %PRODUCTNAME Calc har för dokument kan inte sparas i HTML-format.  
Arkiv - Öppna  
Arkiv - Spara som  
Mata in tal med inledande nollor  
Det finns följande möjligheter om du vill mata in heltal med inledande nollor:  
Mata in talen som text.  
Det är enklast om du matar in talet med ett inledande apostroftecken (t.ex. '0987).  
Apostroftecknet övertas inte i cellen och talet formateras som text.  
Du kan dock inte räkna med det utan vidare.  
Du formaterar cellen med ett talformat som kan se ut så här: \0000.  
Det här formatet (mata in under Format - Cell, i fältet Formatbeskrivning under fliken Tal) definierar visningen i den här cellen som "alltid en nolla först och sedan heltalet, minst tresiffrigt, fyllt med nollor från vänster ".  
Om du i stället t.ex. har importerat en hel kolumn med tal i "textformat", alltså i form av "000123", och nu vill göra "riktiga" tal av dem igen utan inledande nollor i form av "123 ", gör du så här:  
Markera kolumnen där talen i "textformat" står.  
Sätt kolumnens cellformat till "tal"  
Välj Redigera - Sök och ersätt  
I fältet Sök efter matar du in: ^[ 0-9]  
Vid Ersätt med matar du in: &  
Markera Reguljärt uttryck  
Markera Bara markering  
Klicka på Ersätt alla.  
Fixera rader eller kolumner som överskrift  
Gör så här:  
Placera markören i cell A3.  
Välj Fönster - Fixera.  
Om du vill upphäva fixeringen väljer du kommandot igen.  
Fixeringen sker vid det vänstra övre hörnet i den aktuella cellen.  
Om det definierade området inte ska gå att rulla använder du kommandot Fönster - Dela.  
Om du vill skriva ut en viss rad på alla sidor i ett dokument använder du kommandot Format - Utskriftsområden - Redigera.  
Fönster - Fixera  
Fönster - Dela  
Format - Utskriftsområden - Redigera  
Anvisningar för %PRODUCTNAME Calc  
Formatera tabeller och celler  
Mata in värden och formler  
Mata in referenser  
Databasområden i tabeller  
Utvärdering med datapilot o.s.v.  
Skriva ut och förhandsgranskning  
Import och export av dokument  
Övrigt  
Markera flera celler  
Markera rektangulärt område  
Håll ner musknappen och dra från ett hörn till det diagonalt motstående hörnet i området.  
Markera en enskild cell  
Håll ner musknappen och rita upp ett område över två celler, släpp inte musknappen och dra tillbaka till den första cellen igen.  
Nu kan du t.ex. flytta den enskilda cellen med dra-och-släpp.  
Markera flera utspridda celler  
Håll ner Kommando Ctrl -tangenten och klicka på cellerna en och en.  
Förutsättningen är att minst en cell redan har markerats.  
Byta markeringsläge  
På statuslisten kan du byta markeringsläge i fältet som heter STD / UTV / TLF:  
Fältinnehåll  
Effekt vid musklick  
STD  
Cellen markeras om du klickar på den med musen.  
En markering upphävs.  
UTV  
Ett rektangulärt område markeras från den aktuella cellen till cellen som du klickar på när du klickar med musen.  
TLF  
Varje gång du klickar på en cell markeras den och de andra cellerna som du redan har markerat förblir markerade.  
Om du klickar med musen i en markerad cell avmarkeras den.  
Statuslist  
Mata in matrisformel  
Vi visar med hjälp av ett exempel hur du kan mata in en matrisformel, utan att gå in på matrisfunktionernas betydelse.  
Tänk dig att du i kolumnerna A och B har vardera 10 tal under varandra (A1:A10 och B1:B10), och i kolumn C vill du räkna ut summan av de båda talen från samma rad.  
Markera resultatområdet C1:C10.  
Tryck på F2 eller klicka på formellistens inmatningsrad.  
Skriv ett likhetstecken (=).  
Markera de första summandernas område A1:A10.  
Tryck på plustangenten (+).  
Markera de andra summandernas område B1:B10.  
Skift + Kommando Ctrl +Retur.  
Matrisområdet är automatiskt skyddat mot ändringar av innehållet, som radering av rader eller kolumner.  
Men du kan redigera formateringen, t.ex. cellbakgrunden.  
Använda multipel räkneoperation  
Multipla räkneoperationer i kolumner eller på rader  
Om data i dataområdet är placerade under varandra (för kolumner) resp. bredvid varandra (för rader), markerar du dataområdet tillsammans med cellen bredvid eller nedanför som målområde.  
Mata in cellreferensen till den första cellen i dataområdet i fältet Kolumn / Rad.  
I fältet Formler matar du in cellreferensen till formelcellen som refererar till dataområdet.  
Exempel  
Du producerar kramdjur som du säljer för 10 €styck.  
Hur stor vinst gör du per år om du säljer hur många kramdjur?  
Titta på följande tabell:  
A  
B  
C  
D  
E  
F  
1  
Försäljningspris  
10  
Årsförsäljning  
Årsvinst  
2  
Kostnad / styck  
2  
500  
-6000  
3  
Fasta kostnader  
100 000  
1000  
-2000  
4  
Antal  
2000  
1500  
2000  
5  
Vinst  
= B4*( B1 - B2) - B3  
2000  
6000  
Beräkning med en formel och en variabel  
För att beräkna vinsten anger du först ett valfritt tal som antal (antal sålda), i det här exemplet 2000.  
Vinsten räknas ut med formeln Vinst=antal * (försäljningspris - styckkostnader) - fasta kostnader.  
Den här formeln skriver du i B5.  
Ange några försäljningstal i kolumn D, t.ex. i 500-steg från 500 till 5000.  
Markera området D2:E11, alltså värden i kolumn D och de tomma cellerna bredvid i kolumn E.  
Öppna dialogrutan Data - Multipla operationer.  
Med markören i fältet Formler klickar du i cell B5.  
Sätt markören i fältet Kolumn och klicka i cell B4.  
Det betyder:  
B4, antalet, är formelns variabel som ersätts av de markerade kolumnvärdena.  
Stäng dialogrutan med OK.  
Vinsterna visas i kolumn E.  
Beräkning med flera formler samtidigt  
Radera kolumn E.  
Mata in följande formel i C5: = B5 / B4.  
Du beräknar årsvinsten per sålt styck.  
Markera området D2:F11, d.v.s. tre kolumner.  
Öppna dialogrutan Data - Multipla operationer.  
Placera markören i fältet Formler och markera cellerna B5 till C5.  
Sätt markören i fältet Kolumn och klicka i cellen B4.  
Stäng dialogrutan med OK.  
Årsvinsterna visas i kolumn E och årsvinsten per styck i kolumn F.  
Multipel operation via kolumner och rader  
I %PRODUCTNAME kan du utföra multipla räkneoperationer för rader och kolumner tillsammans i s.k. korstabeller.  
Formelcellen ska då hänvisa till det dataområde som ordnats i både rader och kolumner.  
Markera det område som avgränsats genom de båda dataområdena och öppna dialogrutan för multipla räkneoperationer.  
Ange referensen till den första cellen i det område som ordnats radvis i fältet Rad.  
Ange referensen till den första cellen i det område som ordnats kolumnvis i fältet Kolumn.  
Beräkning med två variabler  
Titta på kolumnerna A och B i exempeltabellen ovan.  
Nu ska du inte bara variera kvantiteten i årsproduktionen, utan även försäljningspriset med tanke på vinsten.  
Utöka tabellen som visas ovan.  
I D2 till D11 står talen 500, 1000, o.s.v. till 5000.  
I E1 till H1 skriver du in talen 8, 10, 15, 20.  
A  
B  
C  
D  
E  
F  
1  
Försäljningspris  
10  
8  
10  
2  
Kostnad / styck  
2  
500  
-7000  
-6000  
3  
Fasta kostnader  
10000  
1000  
-4000  
-2000  
4  
Antal  
2000  
1500  
-1000  
2000  
5  
Vinst  
= B4*( B1 - B2) - B3  
2000  
2000  
6000  
Markera området D1:H11.  
Öppna dialogrutan Data - Multipla operationer.  
Placera markören i fältet Formler och klicka i cellen B5.  
Sätt markören i fältet Rad och klicka i B1.  
Det betyder:  
B1, försäljningspriset, är den horisontellt angivna variabeln (med värdena 8, 10, 15 och 20).  
Sätt markören i fältet Kolumn och klicka i cellen B4.  
Det betyder:  
B4, antalet, är den vertikalt angivna variabeln.  
Stäng dialogrutan med OK.  
Vinsterna visas i området E2:H11.  
Eventuellt måste du först trycka på F9 för att uppdatera tabellen.  
Multipla operationer  
Visning av flera tabeller  
Med kommandoknapparna för navigation bläddrar du bland registerflikarna för alla tabeller.  
Om du klickar på kommandoknappen längst till höger i den här gruppen förskjuts visningen av flikar så att du kan se namnet på den sista tabellen.  
För att visa själva tabellen klickar du på namnet på tabellen.  
Om platsen inte räcker till i fönsterkanten för att visa tabellflikarna, kan du förstora den.  
Du gör det genom att dela upp den tillgängliga platsen mellan tabellflikar och horisontell rullningslist.  
Peka på strecket mellan rullningslist och tabellflikar, tryck på musknappen och dra med nertryckt musknapp åt höger.  
Använda flera tabeller  
I förinställningen visar %PRODUCTNAME tre tabeller, "Tabell1" till "Tabell3 ", i alla nya tabelldokument.  
Infoga tabeller  
I snabbmenyn hittar du kommandot Infoga, som används för att infoga en ny tom tabell eller en befintlig tabell från en annan fil framför den aktuella tabellen.  
Markera flera tabeller  
Fliken för den aktuella tabellen visas alltid i vit färg framför de andra flikarna.  
De andra flikarna är grå om de andra tabellerna inte är markerade.  
Du kan markera fler tabeller genom att klicka på deras flikar och samtidigt hålla ner Kommando Ctrl -tangenten.  
Upphäva markering  
Du avmarkerar en tabell genom att klicka på dess flik igen, samtidigt som du håller ner Kommando Ctrl -tangenten.  
Markeringen av den aktuella och synliga tabellen kan inte upphävas.  
Skriva värden i flera tabeller samtidigt  
Om flera tabeller är markerade överförs alla värden som du skriver in i den aktuella tabellen även till de andra markerade tabellerna.  
Det som du matar in i cell A1 i Tabell1 visas alltså även i samma cell i Tabell2, om båda tabellerna är markerade.  
Beräkna funktion över många tabeller (t.ex. medelvärdet av cell A1 över alla tabeller).  
Ange formeln på följande sätt: =MEDEL( tabell1.A1:tabell50.A1).  
Nu bildas medelvärdet i formelcellen för alla A1-celler i dina 50 tabeller.  
Infoga och redigera anteckningar  
Varje cell kan innehålla en anteckning som du infogar via menypunkten Infoga - Anteckning.  
En liten röd kvadrat indikerar att cellen innehåller en anteckning.  
Anteckningen visas när du pekar med musen på cellen, under förutsättning att du har aktiverat Tips eller Aktiv hjälp på menyn Hjälp.  
Om du markerar cellen kan du välja Visa anteckning på cellens snabbmeny.  
Då visas anteckningen hela tiden tills du upphäver kommandot Visa anteckning på cellens snabbmeny.  
Du redigerar en anteckning som alltid visas genom att klicka i den.  
Om du raderar hela anteckningstexten raderas anteckningen.  
Du kan också radera en anteckning i dialogrutan Redigera - Radera innehåll som du öppnar med tangenten Delete.  
Du kan visa och dölja anteckningsmarkören under Verktyg - Alternativ - Tabelldokument - Vy.  
Infoga - Anteckning  
Skriva ut tabelldetaljer  
När du skriver ut en tabell kan du välja vilka detaljer som ska skrivas ut:  
Radhuvuden och kolumnhuvuden  
Tabellgitter  
Anteckningar  
Objekt och grafik  
Diagram  
Ritobjekt  
Formler  
Gör så här för att välja detaljer:  
Växla till tabellen som du vill skriva ut.  
Välj Format - Sida.  
Kommandot visas inte om tabellen är skrivskyddad.  
Klicka då först på ikonen Redigera fil på funktionslisten.  
Klicka på fliken Tabell.  
Välj detaljerna som ska skrivas ut i området Skriv ut och klicka på OK.  
Skriv ut dokumentet.  
Visa - Förhandsvisning av sidbrytningar  
Definiera antal utskriftssidor  
%PRODUCTNAME Calc kommer att skriva ut den aktuella tabellen jämt fördelad på flera sidor om den är för stor för en enda utskriftssida.  
Eftersom den automatiska sidbrytningen inte alltid sker på det ställe som du skulle ha valt, kan du även definiera uppdelningen av sidor själv:  
Växla till tabellen som ska skrivas ut.  
Välj Visa - Förhandsvisning av sidbrytningar.  
Du ser den automatiska uppdelningen av tabellen på utskriftssidor.  
Utskriftsområdena som har skapats automatiskt är markerade med blåa linjer, utskriftsområden som har definierats av användaren med ljusblå linjer.  
Sidbrytningarna (radbrytningar och kolumnbrytningar) markeras med svarta linjer.  
Du kan flytta de blåa linjerna med musen.  
På snabbmenyn finns det fler möjligheter, bl.a. att lägga till ett ytterligare utskriftsområde, upphäva utskriftsområden, upphhäva skalning och infoga fler manuella rad - och sidbrytningar.  
Visa - Förhandsvisning av sidbrytningar  
Skriva ut tabell i liggande format  
När du ska skriva ut en tabell har du många interaktiva möjligheter om du väljer Visa - Förhandsvisning av sidbrytning.  
Om du vill skriva ut tabellen på papper i liggande format, gör du så här:  
Växla till tabellen som du vill skriva ut.  
Välj Format - Sida.  
Kommandot visas inte om tabellen är skrivskyddad.  
Klicka då först på ikonen Redigera fil på funktionslisten.  
Klicka på fliken Sida.  
Välj pappersformatet Liggande och klicka på OK.  
Välj Arkiv - Skriv ut.  
Dialogrutan Skriv ut öppnas.  
Allt efter skrivardrivrutin och operativsystem kan du behöva klicka på kommandoknappen Egenskaper och ställa om din skrivare till liggande format.  
Välj vilka sidor som ska skrivas ut under Utskriftsområde i dialogrutan Skriv ut:  
Allt - alla tabeller skrivs ut.  
Sidor - du anger sidorna som ska skrivas ut.  
Sidorna räknas alltid från den första tabellen.  
Om du ser i förhandsvisningen av sidbrytningar att Tabell1 skrivs ut på 4 sidor, och du vill skriva ut de första båda sidorna av Tabell2, anger du 5-6 här.  
Markering - bara markeringen skrivs ut.  
Om celler är markerade skrivs de ut.  
Om inga celler är markerade, skrivs alla tabeller ut vars namn är markerade (på tabellflikarna).  
Du ändrar markeringen genom att hålla ner Ctrl-tangenten och klicka på ett av tabellnamnen.  
Om du har definierat ett eller flera utskriftsområden under Format - Utskriftsområden, skrivs bara innehållet i de här utskriftsområdena ut.  
Visa - Förhandsvisning av sidbrytningar  
Skriva ut rad eller kolumn på varje sida  
Du har en tabell som skrivs ut på fyra sidor på grund av sin omfattning.  
Utskriftssidorna är ordnade på följande sätt:  
Sida 1  
Sida 3  
Sida 2  
Sida 4  
De båda översta raderna i tabellen ska inte bara skrivas ut på sidan 1 och 3 utan även som översta rader på sidan 2 och 4.  
Den första kolumnen A ska inte bara skrivas ut på sidan 1 och 2 utan även på sidan 3 och 4.  
Välj Format - Utskriftsområden - Redigera.  
Dialogrutan Redigera utskriftsområden öppnas.  
Klicka på ikonen längst till höger i området Upprepningsrad.  
Dialogrutan förminskas så att du kan se mer av tabellen.  
Markera de två första raderna genom att t.ex. klicka i cell A1 och dra till A2.  
I den förminskade dialogrutan står $1:$2.  
Raderna 1 och 2 är nu upprepningsrader.  
Klicka på ikonen längst till höger i området Upprepningsrad.  
Dialogrutan förstoras.  
Om du även vill ha kolumnen A som upprepningskolumn, klickar du på ikonen längst till höger i området Upprepningskolumn.  
Klicka i kolumn A (inte på kolumnhuvudet).  
Klicka på ikonen längst till höger i området Upprepningskolumn igen och sedan på OK.  
Upprepningsrader är rader från tabellen.  
Sidhuvuden och sidfötter som skrivs ut på alla sidor kan du definiera oberoende av dem via Format - Sida.  
Visa - Förhandsvisning av sidbrytningar  
Format - Utskriftsområden - Redigera  
Format - Sida - (Sidhuvud / Sidfot)  
Adresser och referenser, absoluta och relativa  
Relativ adressering  
Med A1 adresseras cellen i kolumn A och rad 1.  
Ange slutligen den högra undre cellen av området.  
Det kvadratiska området av de första fyra cellerna i hörnet uppe till vänster heter då A1:B2.  
Vid den här typen av adressering av ett område är referensen till A1:B2 en relativ referens.  
Relativ betyder här att referensen till det här området anpassas när du kopierar formlerna.  
Absolut adressering  
I motsats till relativ adressering finns den absoluta referensen som skrivs på följande sätt: $A$1:$B$2.  
Det står alltså ett dollartecken framför varje angivelse som skall användas absolut.  
Om du trycker på Skift+F4 kan %PRODUCTNAME skriva om den aktuella referensen där markören står i inmatningsraden från relativ till absolut och tillbaka.  
Om du inleder med en relativ adress som A1, gäller följande:  
Första gången du trycker sätts rad och kolumn till absolut ($A$1), nästa gång du trycker bara raden (A$1), sedan bara kolumnen ($A1) och sedan blir referensen relativ i båda riktningar igen (A1).  
%PRODUCTNAME Calc visar referenserna till en formel.  
Om du t.ex. klickar på formeln =SUMMA( A1:C5;D15:D24) i en cell, markeras de båda referensområdena i tabellen i färg.  
Formeldelen "A1:C5" kan till exempel visas i blått och det aktuella cellområdet är inramat med samma blåton.  
Nästa formeldel "D15:D24" kan vara markerad på samma sätt i rött.  
När används relativa och när används absoluta referenser?  
Vad utmärker en relativ referens?  
Vi antar att du vill beräkna summan av cellerna i området A1:B2 i cell E1.  
Formeln som du matar in i E1 skulle alltså vara =SUMMA( A1:B2).  
Nu bestämmer du dig senare för att infoga en kolumn till framför kolumn A.  
Elementen som du vill summera, står sedan plötsligt i B1:C2 och formeln står inte längre i E1, utan i F1.  
Du måste alltså kontrollera och korrigera alla formler i tabellen - och eventuellt i andra tabeller - när du har infogat den nya kolumnen.  
Som tur är gör %PRODUCTNAME det här arbetet åt dig när rader infogas och raderas.  
Formeln =SUMMA( A1:B2) korrigeras automatiskt till =SUMMA(B1:C2) om en ny kolumn A har infogats.  
De absoluta och relativa referenserna anpassas alltid automatiskt i %PRODUCTNAME Calc när referensdataområdet förskjuts.  
Men du måste se upp när du kopierar formler: då anpassas nämligen bara de relativa referenserna och inte de absoluta.  
Absoluta referenser sätter du in när beräkningar refererar till exakt en cell i din tabell där t.ex. ett procentvärde står.  
Om en formel, som refererar till just den här cellen, kopieras relativt neråt, förskjuts referensen också neråt om du inte har satt cellkoordinatorerna absolut.  
Förutom när nya rader och kolumner infogas, kan referenser också ändras när du har matat in en formel som refererar till bestämda celler och sedan kopierar den här formeln för ett annat område i tabellen.  
Tänk dig att du har matat in summan av de ovanstående cellerna i formeln =SUMMA( A1:A9) på rad 10.  
Om du nu också vill beräkna summorna i kolumnerna som står bredvid till höger, kan du helt enkelt kopiera den här formeln åt höger.  
För kopian av formeln som står i kolumn B, hittar du sedan den automatiskt korrigerade formeln =SUMMA( B1:B9).  
Byta namn på en tabell  
Klicka på tabellnamnet som du vill ändra, t.ex. på "Tabell1".  
Öppna snabbmenyn och välj Byt namn.  
Du ser en dialogruta där du kan mata in ett nytt namn för tabellen.  
Mata in det nya namnet på tabellen och klicka på OK.  
Alternativt kan du också hålla ner Alternativtangenten Alt-tangenten och klicka på ett tabellnamn och sedan mata in det nya namnet direkt.  
Det får innehålla mellanslag.  
Namnet på en tabell är inte beroende av namnet på tabelldokumentet.  
Dokumentet kan innehålla upp till 256 enskilda tabeller som har olika namn.  
Använda avrundade tal  
I %PRODUCTNAME Calc visas alla decimaltal avrundade till två decimaler.  
Går det att ändra för markerade celler?  
Markera alla celler vars talformat du vill ändra.  
Välj Format - Cell och klicka på fliken Tal.  
Välj Tal i fältet Kategori.  
Ändra Antal decimaler under Alternativ och avsluta dialogrutan med OK.  
Går det att ändra en gång för alla?  
Välj Verktyg - Alternativ - Tabelldokument.  
Klicka på fliken Beräkna.  
Ändra Antal decimaler och avsluta dialogrutan med OK.  
Går det att räkna med de visade avrundade värdena i stället för de interna exakta värdena?  
Välj Verktyg - Alternativ - Tabelldokument.  
Klicka på Beräkna.  
Markera rutan Precision som visat och avsluta dialogrutan med OK.  
Fliken tal  
Beräkna  
Ändra radhöjd eller kolumnbredd  
Du kan ändra radhöjden med musen eller i en dialogruta.  
Det som beskrivs här för rader och radhöjd gäller även för kolumner och kolumnbredd.  
Ändra radhöjd eller kolumnbredd med musen  
Klicka på strecket nedanför den aktuella raden i området med radhuvuden, håll ner musknappen och dra nedåt eller uppåt så ändras radhöjden.  
Den optimala radhöjden väljer du genom att dubbelklicka på strecket nedanför raden.  
Ändra radhöjd eller kolumnbredd i dialogruta  
Klicka på raden så att den fokuseras.  
Öppna snabbmenyn på radhuvudet i den vänstra kanten.  
Du ser bl.a. kommandona Radhöjd och Optimal radhöjd som öppnar en dialogruta.  
Radhöjd  
Optimal radhöjd  
Kolumnbredd  
Optimal kolumnbredd  
Använda scenarion  
Scenarion är viktiga hjälpmedel för att se siffror som är beroende av varandra och beräkningarna som de resulterar i.  
Ändra vissa grundläggande förutsättningar i tabellen och titta på det nya resultatet.  
Du kan ge scenariot som du har skapat ett namn och sedan jämföra det med andra scenarion.  
Använda färdiga scenarion  
Det finns ett utarbetat exempel med scenarion.  
Välj Arkiv - Nytt - Mallar och dokument och klicka där på Exempel.  
Öppna tabellexemplen.  
Du ser nu de medföljande tabelldokumenten.  
Dubbelklicka på dokumentet med Recar i namnet.  
Du ser nu en exempeltabell där redan flera scenarion har skapats.  
Områdena där de olika utgångsvärdena beroende på scenario står, är inramade.  
Du väljer ut respektive giltigt scenario i listrutan som finns i övre kanten på varje ram.  
Alternativt kan du välja ut scenarierna i Navigator:  
Öppna Navigator, t.ex. med tangenten F5 eller med ikonen Navigator på funktionslisten.  
I Navigator klickar du på ikonen Scenarion (ikonen med utrops - och frågetecken).  
Du ser nu de definierade scenarierna i Navigator med kommentarerna som fördes in där när scenarierna skapades.  
Skapa egna scenarion  
För att skapa ett scenario måste du markera alla celler som innehåller data för scenariot.  
I vårt exempel kan du skapa ett ytterligare scenario som t.ex. heter "Hög dollarkurs".  
Gör så här:  
Markera alla dataceller som redan framhävs av det bestående scenariots ram.  
Om uppgifterna inte finns i ett genomgående område, utan är fördelade över tabellen, kan du även göra en multimarkering.  
Det gör du genom att hålla ner Kommando Ctrl -tangenten medan du klickar på cellerna.  
Men i vårt exempel behöver du bara markera området F18:F23.  
Du ser dialogrutan Skapa scenario.  
Stäng dialogrutan med OK.  
Ditt nya scenario är automatiskt aktiverat.  
Ändra värdena i ramarna till värdena som skall gälla för ditt nya scenario.  
Ändra i det här fallet dollarkursen och alla värden som enligt din mening kan påverkas av den, t.ex. ekonomisk tillväxt och försäljningspriser.  
Du ser genast effekterna på siffrorna.  
Spår till efterträdaren.  
Om du vill veta vilka värden som påverkar vilka andra värden i scenarierna, väljer du Verktyg - Detektiv - Spår till efterträdaren.  
Du ser sedan pilar till cellerna som är direkt beroende av den aktuella cellen.  
Skapa scenarion  
Använda sorteringslistor  
Mata in texten "jan" eller "januari "i en tom tabellcell.  
Dra i högra hörnet på ramen runt cellen åt höger eller neråt över flera celler.  
När du släpper musknappen fylls de överstrukna cellerna med den definierade serien av månadernas namn.  
Här kan du även mata in egna sorteringslistor, till exempel en lista över ditt företags filialer.  
Om du behöver den här listan senare, t.ex. som tabellrubriker, räcker det att mata in det första namnet och utöka inmatningen genom att dra med musen.  
Sorteringslistor  
Filter: använda specialfilter  
Kopiera överskrifterna i det tabellområde som ska filtreras till en tom plats i tabellen och ange kriterierna nedanför dem.  
Data som står horisontellt bredvid varandra kombineras då alltid logiskt med OCH, och data som står vertikalt under varandra kombineras alltid logiskt med ELLER.  
Om du har skapat en sådan filtermatris markerar du tabellområdet som ska filtreras, öppnar Specialfilter-dialogrutan och väljer sedan definitionen av specialfiltret.  
Sedan klickar du på OK och ser då att bara de rader i ursprungstabellen visas, vars innehåll stämde med sökkriterierna.  
Alla andra rader är dolda och kan visas igen med kommandot Format - Rad - Visa.  
Exempel  
Ladda ett tabelldokument med så många dataposter som möjligt.  
Vi utgår här från ett fiktivt dokument, Omsättning, men du kan lika gärna använda vilket annat dokument som helst.  
Dokumentet ser ut ungefär så här:  
A  
B  
C  
D  
E  
1  
Månad  
Standard  
Business  
Lyx  
Suite  
2  
januari  
12560  
200500  
24000  
17000  
3  
februari  
16000  
180300  
36200  
22000  
4  
mars  
17000  
och så vidare...  
Kopiera rad 1 med överskrifterna = datafältnamnen till rad 20, till exempel.  
Ange filtervillkoren som är länkade med ELLER på rad 21, 22 och så vidare.  
Området skulle kunna se ut så här:  
A  
B  
C  
D  
E  
20  
Månad  
Standard  
Business  
Lyx  
Suite  
21  
=" januari "  
22  
<160000  
Här definierar du att bara de rader ska visas som antingen har värdet "januari" i fältet Månad ELLER ett värde under 160000 i fältet Standard.  
Välj kommandot Data - Filter - Specialfilter och markera sedan området A20:E22 med hjälp av musen.  
Nu visas bara de filtrerade raderna i tabellområdet.  
De andra raderna döljs.  
Filter: använda standardfilter  
Med hjälp av posten - Standard - i AutoFilter eller med kommandot Data - Filter - Standardfilter öppnar du dialogrutan Standardfilter.  
Här anger du upp till tre villkor för filtreringen.  
Alternativen i dialogrutan Standardfilter beskrivs utförligt i %PRODUCTNAME -hjälpen.  
I illustrationen har vi definierat att bara de rader i det markerade området ska visas, där datafältet "Månad" har värdet "januari "och samtidigt datafältet "Standard" har ett värde som är större eller lika med 160000.  
Data - Filter - Standardfilter  
Upphöjd / nedsänkt text  
Markera tecknen som ska vara upphöjda eller nedsänkta.  
Om du t.ex. vill skriva H2O markerar du 2:an i cellen (inte på inmatningsraden).  
Öppna snabbmenyn till de markerade tecknen och välj kommandot Tecken.  
Dialogrutan Tecken öppnas.  
Klicka på fliken Teckenposition.  
Välj alternativet Nedsänkt och klicka på OK.  
Snabbmeny - Tecken - Teckenposition  
Rotera tabell (transponera)  
Finns det ett sätt att "rotera" en tabell i %PRODUCTNAME Calc så att rader blir till kolumner och tvärtom?  
Markera först tabellområdet som du vill transponera.  
Välj meny Redigera - Klipp ut.  
Upphäv markeringen.  
Sätt markören i cellen som skall vara den vänstra övre cellen för resultatet.  
Välj meny Redigera - Klista in innehåll.  
I dialogrutan aktiverar du sedan rutan Klistra in allt i området Urval och rutan Transponera i området Alternativ.  
När du nu klickar på kommandoknappen OK byter kolumner och rader plats med varandra.  
Klistra in innehåll  
Ändra visning av tabell  
Så döljer du kolumn - och radhuvuden i en tabell permanent.  
Välj Verktyg - Alternativ - Tabelldokument, och sedan Vy.  
Bekräfta med OK.  
Så döljer du gitterlinjerna  
Välj Verktyg - Alternativ - Tabelldokument, och sedan Vy.  
Avmarkera Gitterlinjer.  
Bekräfta med OK.  
Formatera tal som text  
Du kan också mata in tal i formatet "Text".  
Formatera ett område av celler med formatet "Text" (snabbmeny Formatera celler - flik Tal, kategori Text) och mata sedan in siffror i de här cellerna, så tolkas de genast som texttecken.  
Det går inte räkna med tal som omvandlats till texttecken!  
Om du redan har matat in normala tal i celler och sätter formatet på cellerna till "Text" i efterhand, förblir talen tal och konverteras alltså inte.  
Det är bara om du matar in nya siffror eller redigerar de redan inmatade talen som de omvandlas till texttecken.  
Om du vill mata in ett tal som texttecken direkt, inleder du inmatningen med apostrof ('), som t.ex. för årsangivelserna i kolumnöverskrifter '1999, '2000 och '2001.  
Apostrofen signalerar att inmatningen ska behandlas som text.  
Den här inmatningen är t.ex. praktisk om du matar in ett telefonnummer eller ett postnummer som börjar med en nolla.  
I normalt talformat skulle det inte vara möjligt att använda inledande nolla.  
Format - Cell - Tal  
Rotera text  
Markera cellerna vars text du vill rotera.  
Välj kommandot Format - Cell.  
Dialogrutan Cellattribut öppnas.  
Klicka på fliken Justering.  
I området Skrivriktning väljer du i vilken riktning texten ska roteras genom att klicka på cirkeln.  
Klicka på OK.  
Om kommandoknappen ABCD är intryckt i området Skrivriktning skrivs texten lodrätt tecken för tecken.  
Format - Cell  
Format - Cell - Justering  
Skriva text på flera rader  
Med tangentkombinationen Kommando Ctrl +Retur infogar du en manuell radbrytning när du skriver.  
Den här tangentkombinationen fungerar bara direkt i cellen, inte på inmatningsraden.  
Om texten ska brytas automatiskt i den högra kanten av cellen gör du så här:  
Markera alla celler där texten ska brytas i den högra kanten.  
Klicka sedan på OK.  
Format - Cell  
Definiera funktion  
Du kan använda användardefinierade funktioner i %PRODUCTNAME Calc på följande sätt:  
I %PRODUCTNAME -hjälpen hittar du information om du vill programmera funktionerna som Add-in.  
Den här metoden förutsätter att du har lite mer erfarenhet av programmering.  
Med hjälp av Basic-IDE:n kan du definiera egna funktioner även om du inte har erfarenhet av programmering.  
Beskrivningen finns på de följande raderna:  
I det här exemplet definierar vi en funktion VOL( a; b; c), som beräknar volymen för en kvader med kantlängderna a, b och c.  
Definiera egen funktion i Basic-IDE  
Välj Verktyg - Makro.  
Dialogrutan Makro öppnas.  
Klicka på kommandoknappen Redigera.  
Du ser Basic-IDE:n.  
Ange funktionen som på bilden.  
Stäng Basic-IDE-fönstret med kommandoknappen på titellisten.  
Din funktion sparas automatiskt i standardmodulen och är sedan alltid tillgänglig i ditt %PRODUCTNAME.  
Om du använder funktionen i ett Calc-dokument som ska användas även på andra datorer, kan du kopiera funktionen till Calc-dokumentet.  
Beskrivningen finns nedan under rubriken "Kopiera egen funktion till ett dokument".  
Använda egen funktion i %PRODUCTNAME Calc  
När du har definierat funktionen VOL( a; b; c) i Basic-IDE:, kan du använda den precis som de installerade funktionerna i %PRODUCTNAME Calc.  
Öppna ett %PRODUCTNAME Calc-dokument och mata t.ex. in några tal i kolumnerna A, B och C.  
Sätt markören i cell D1 och mata in följande:  
=VOL( A1;B1;C1)  
Funktionen utvärderas och du ser resultatet i cell D1.  
Kopiera egen funktion till ett dokument  
I steg 2 till "Definiera egen funktion i Basic-IDE" klickade du på Redigera i dialogrutan Makro.  
Standardmodulen är soffice - Standard - Modul1 som är utvald i fältet Makro från.  
Standardmodulen ligger lokalt i din användarkatalog.  
Om du vill kopiera den egna funktonen till ett Calc-dokument, gör du så här:  
Välj Verktyg - Makro.  
Välj modulen soffice - Standard - Modul1 i fältet Makro från.  
Klicka på Redigera.  
I Basic-IDE:n markerar du källtexten till din egen funktion och kopierar den till urklippet.  
Stäng Basic-IDE:n.  
Välj Verktyg - Makro.  
Välj modulen (Namn på Calc-dokumentet) - Standard - Modul1 i fältet Makro från.  
Klicka på Redigera.  
Klistra in innehållet i urklippet i Basic-IDE:n till dokumentet.  
Byt till "Hjälp till %PRODUCTNAME Basic", sök sedan efter "Integrerad utvecklingsmiljö (IDE)"  
Validitet för cellinnehåll  
Du kan definiera för varje cell i förväg vilken typ av innehåll som ska vara giltigt för den här cellen.  
På så sätt gör du det lättare för användarna att använda tabellen på rätt sätt.  
Giltighetsregeln används när ett nytt värde anges.  
Om det redan finns ett (ogiltigt) värde i cellen eller om du placerar ett värde i cellen genom att dra och släppa eller kopiera och klistra in gäller inte giltighetsregeln.  
Du kan välja Verktyg - Detektiv - Ringa in ogiltiga data för att se om det finns några värden som inte är giltiga.  
Det finns detaljerad information om kommandot Data - Validitet i %PRODUCTNAME -hjälpen.  
Så här arbetar du med giltighet för cellinnehåll  
1.  
Markera de celler för vilka du vill definiera en ny giltighetsregel.  
Du kan också göra en multimarkering genom att klicka på alla önskade celler, samtidigt som du håller ner Kommando Ctrl -tangenten.  
Giltighetsregeln är en del av en cells format.  
Du kan kopiera giltighetsregeln till andra celler med Redigera - Kopiera och Redigera - Klistra in innehåll, urval "Format".  
2.  
Välj Data - Validitet....  
Dialogrutan Validitet visas.  
3.  
Klicka på fliken Kriterier och ange de villkor som värdena i cellen måste uppfylla.  
Redan befintliga värden påverkas inte.  
4.  
I listrutan Tillåt är "Alla värden" förinställning.  
Det innebär att det inte finns några inskränkningar.  
Du kan välja mellan fler möjligheter: heltal, decimal, datum, tid och textlängd.  
5.  
Med detta val anger du det första villkoret.  
Om du väljer "Heltal" är värden som t.ex. "12,5 "inte tillåtna, även om de inte skulle strida mot de övriga villkoren.  
Om du väljer "Datum" är datumangivelser tillåtna både i form av "1.1.00 "och av ett seriellt datumtal.  
Liknande gäller för "Tid", där bara inmatningar av typen "12:00" eller seriella tidstal är tillåtna.  
Med "Textlängd" definierar du att enbart text är tillåtet som cellinnehåll.  
6.  
När du har angett det första villkoret under Tillåt väljer du nästa villkor under Data.  
Beroende på vilket villkor du har valt visar dialogrutan fler textfält som heter Värde, Minimum och Maximum, där du kan specificera villkoret ytterligare.  
7.  
Några tänkbara villkor som kan formuleras under denna flik ser ut så här: "Heltal större än 1", "Decimal mellan 10 och 12,5", "Datum mindre än eller lika med 1.1.2000", "Tid inte lika med 00:00", "Textlängd större än 2 tecken".  
Därmed har du definierat villkoret för de värden som därefter matas in i denna cell.  
Om det skulle förekomma avvikelser visar %PRODUCTNAME ett standardmeddelande.  
Du kan ge användaren mer hjälp genom att fylla i mer information under de båda andra flikarna.  
Under fliken Inmatningshjälp anger du rubriken och texten till den tipshjälp som ska visas när cellen markeras.  
Under fliken Felmeddelande väljer du vad som ska hända vid en felaktig inmatning.  
Det gamla innehållet i cellen bibehålls.  
Om du väljer åtgärden "Varning" eller "Information "öppnas en dialogruta där du kan avbryta inmatningen (cellens gamla värde bibehålls) eller godkänna den (det nya värdet accepteras trots att det strider mot giltighetsregeln).  
Om du väljer åtgärden "Makro" kan du ange ett makro, som utförs vid felaktig inmatning, med hjälp av kommandoknappen Genomsök.  
Om du ändrar åtgärden som är knuten till en cell under fliken Felmeddelande och avslutar dialogrutan med OK måste du först markera en annan cell innan ändringen blir verksam.  
Data - Validitet  
Namnge celler  
Du har t.ex. matat in en aktuell omräkningsfaktor på 2,34 i cell X1.  
Du kan göra formlerna som använder den här faktorn lättare att läsa genom att ge cellen X1 ett namn.  
Formeln lyder då t.ex. inte längre = A1 * X1 utan = A1 * omräkningsfaktor.  
Markera cell X1 (i det här exemplet), sedan väljer du menykommandot Infoga - Namn - Definiera.  
Dialogrutan Definiera namn öppnas.  
Mata till exempel in namnet i textfältet Omräkningsfaktor.  
Klicka på Lägg till och stäng dialogrutan.  
Om du nu börjar mata in namnet Omräkningsfaktor i en formel ser du hela namnet som tipshjälp när du har matat in de första tecknen.  
Tryck på returtangenten om du vill använda namnet från tipshjälpen.  
Om flera namn börjar med samma tecken kan du bläddra igenom alla namnen med tabbtangenten.  
Infoga - Namn - Definiera  
Infoga externa data i tabell  
Med hjälp av importfiltret Webbsidessökning i kategorin %PRODUCTNAME Calc-filter infogar du tabeller från HTML-dokument i ett %PRODUCTNAME Calc-tabelldokument.  
Du kan även använda samma metod när du ska infoga områden som är definierade med namn från ett %PRODUCTNAME Calc-tabelldokument.  
Det finns följande infogningsmetoder:  
Infoga via dialogruta  
Placera cellmarkören i cellen från vilken du vill infoga det nya innehållet.  
Välj Infoga - Externa data.  
Dialogrutan Externa data öppnas.  
Ange HTML-dokumentets URL eller namnet på tabelldokumentet i kombinationsfältet.  
Du kan välja fil med hjälp av en dialogruta.  
Den valda filen laddas i bakgrunden (osynlig).  
Sedan kan du välja områdena eller tabellerna från filen i den stora listrutan i dialogrutan.  
Om du vill definierar du att områdena eller tabellerna ska uppdateras var n sekund.  
Infoga med Navigator  
1.  
Öppna två dokument: %PRODUCTNAME Calc-tabelldokumentet där du vill infoga externa data (måldokument) och dokumentet från vilket externa data ska hämtas (källdokument).  
2.  
Öppna Navigator i måldokumentet.  
3.  
I det undre kombinationsfältet i Navigator väljer du ut källdokumentet.  
Navigator visar nu områdesnamnen och databasområdena resp. tabellerna som finns i källdokumentet.  
4.  
Välj draläget Infoga som länk i Navigator.  
5.  
Dra de externa data som du vill använda från Navigator till måldokumentet.  
Om du har laddat ett HTML-dokument med filtret Webbsidessökning som källdokument, finns tabellerna i Navigator, kallade för "HTML_table1" o.s.v. och dessutom två områdesnamn som har skapats:  
HTML_all - betecknar hela dokumentet  
HTML_tables - betecknar alla HTML-tabeller i dokumentet  
Redigera externa data  
Öppna dialogrutan Redigera - Länkar.  
Här kan du redigera länken till externa data.  
Dialogrutan Externa data  
Årtal 19xx / 20xx  
Årtal i datumangivelser anges ofta med två siffror.  
Internt administreras årtalen med fyra siffror av %PRODUCTNAME så att resultatet vid beräkningen av differensen mellan 99-01-01 och 01-01-01 blir rätt, d.v.s. två år.  
Under Verktyg - Alternativ - %PRODUCTNAME - Allmänt kan du ställa in till vilket år ett tvåsiffrigt årtal "xx" ska visas som "20xx ".  
Det betyder att om du anger datumet 30-01-01. eller högre, behandlas det internt som 1930-01-01 eller högre.  
Alla mindre årtal gäller i följande århundrade, 20-01-01 omvandlas t.ex. till 2020-01-01.  
Välkommen till %PRODUCTNAME Calc-hjälpen  
Hjälp till %PRODUCTNAME Calc  
Lista över kategorier och funktioner  
Hjälp till hjälpen  
Menyer  
När du arbetar med tabelldokument finns kommandon som används till att redigera dokumenten på menylisten.  
Arkiv  
På den här menyn finns kommandon som används till att hantera dokument i sin helhet.  
Du kan t.ex. skapa ett nytt dokument, öppna, stänga och skriva ut dokument, ange dokumentegenskaper med mera.  
När Du vill avsluta %PRODUCTNAME klickar du på menykommandot Avsluta.  
Öppna  
Spara som  
Versioner  
Egenskaper  
Skriv ut  
Skrivarinställning  
Redigera  
Här finns även olika funktioner för att redigera förteckningar och integrerade objekt.  
Dessutom hittar du här kommandon för att fylla i celler automatiskt, radera innehåll, celler och tabeller och flytta och kopiera tabeller.  
Klistra in innehåll...  
Jämför dokument...  
Sök och ersätt...  
Sidhuvud och sidfot...  
Radera innehåll...  
Radera celler...  
Radera tabell...  
Kopiera / Flytta tabell...  
Länkar...  
Image map  
Visa  
Visa-menyn innehåller kommandon som används till att styra hur tabelldokumentfönstret och dokumentinnehållet ser ut på bildskärmen.  
Här kan du bestämma vilka av symbollisterna som ska visas eller i vilken skala dokumentet ska visas.  
Skala...  
Infoga  
På den här menyn finns alla kommandon som används till att infoga nya element i dokumentet, som t.ex. celler, rader, kolumner, tabeller och namn på celler, samt en lista över kategorier och funktioner.  
Du kan även infoga specialtecken, grafik, objekt från andra tillämpningar o.s.v. här.  
Celler...  
Tabell...  
Specialtecken...  
Hyperlänk  
Funktion...  
Funktionslista  
Anteckning Anteckning...  
Diagram...  
Ram  
Format  
På menyn Format finns kommandon som du behöver till att formatera det för tillfället markerade objektet i dokumentet.  
Vilka menykommandon som visas beror på vilket objekt som är markerat.  
Om det aktuella objektet är en ram eller en grafik, så visar menyn kommandona som behövs för detta objekt.  
Dessutom innehåller menyn funktioner som används till att hantera formatmallar, t.ex. mallkatalogen och Stylist.  
Cell...  
Linje...  
Yta...  
Text...  
Position och storlek...  
Kontrollfält...  
Formulär...  
Tecken...  
Stycke...  
Sida...  
Mallkatalog...  
AutoFormat...  
Villkorlig formatering...  
Verktyg  
Här startar du rättstavningskontrollen för de texter som finns i cellerna eller öppnar synonymordlistan som ger dig förslag på alternativa ord.  
Här kan du även använda Detektiv-funktionen för att leta efter tabellreferenser och fel och starta målvärdessökningen eller definiera scenarion.  
Dessutom kan du starta makro-programmeringen här och göra inställningar för symbollister, menyer och tangentbordet och allmänna förinställningar för programmet.  
Synonymordlista...  
Målvärdessökning...  
AutoKorrigering...  
Målvärdessökning  
Scenarion...  
Datakällor  
Makro...  
Anpassa...  
Fönster  
På Fönster-menyn hittar du kommandon som används till att öppna, dela och fixera fönster.  
Data  
Här hittar du kommandona för att redigera data i tabelldokument.  
Här kan du bl.a. definiera områden, sortera och filtrera data, beräkna resultat, disponera data och starta datapiloten.  
Definiera område...  
Välj område...  
Sortera...  
Delresultat...  
Validitet...  
Multipla räkneoperationer...  
Konsolidera...  
Uppdatera område...  
Symbollister  
Här hittar du en beskrivning av elementen som finns på symbollisterna i ett aktivt tabelldokument.  
Tabellobjektlist  
Tabellobjektlisten innehåller de vanligaste funktionerna för direkt teckenformatering, d.v.s. formatering utan användning av formatmallar, i tabelldokument.  
Med kommandot Format - Standard kan du ta bort alla direkta formateringar i de markerade cellerna.  
Teckenfärg  
Vänsterjusterad  
Justering centrerat horisontellt  
Högerjusterad  
Marginaljusterad  
Justera överkant  
Justera centrerat vertikalt  
Justera nederkant  
Objektlisten för ett markerat objekt  
Objektlisten för markerade objekt innehåller de funktioner som är viktigast för att du ska kunna formatera och justera dessa objekt.  
Den här objektlisten visas om du har markerat ett objekt i tabellen, ett grafiskt objekt eller en teckning.  
Du kan konfigurera den och lägga till och ta bort så många ikoner som du vill om du väljer menykommandot Visa - Symbollister - Redigera....  
Samma dialogruta öppnar du med Verktyg - Anpassa... och kommandoknappen Redigera... under fliken Symbollister.  
Linjestil  
Linjebredd  
Linjefärg  
Ytstil / -fyllning  
Objektlisten med textmarkören i ett objekt  
Om textmarkören t.ex. står i en infogad textram, visas ikonerna för textformatering på denna objektlist.  
Den här objektlisten visas även om du sätter textmarkören i ett objekt genom att dubbelklicka när du vill skriva text i objektet.  
Teckensnittsfärg  
Radavstånd:  
1  
Radavstånd:  
1,5  
Radavstånd:  
2  
Vänsterjusterad  
Centrerad  
Högerjusterad  
Marginaljustering  
Upphöjt  
Nedsänkt  
Teckenattribut  
Format: stycke  
Formellist  
Formellisten använder du när du ska mata in matematiska formler.  
Statuslist  
Statuslisten visar information om det aktuella dokumentet och innehåller några kommandoknappar med specialfunktioner.  
Du kan konfigurera statuslisten (under Verktyg - Anpassa...) på samma sätt som övriga lister.  
Normalt visas fält som har följande betydelse:  
Förhandsgranskningslist  
Förhandsgranskningslisten visas när du har aktiverat förhandsgranskningen för det aktuella dokumentet (via kommandot Förhandsgranskning på menyn Arkiv).  
Sidformat  
Grafikobjektlisten  
Om ett grafikobjekt är markerat i ett dokument visas grafikobjektlisten.  
Verktygslist  
Här har du tillgång till de viktigaste funktionerna.  
Formulär  
Temaurval  
Sökning på / av  
Sortera  
Funktioner i %PRODUCTNAME Calc  
Här får du en kort överblick över några viktiga funktioner i %PRODUCTNAME Calc.  
Räkna  
Det har tabeller i vars celler du kan mata in texter, tal och formler och genomföra enkla och komplexa beräkningar.  
Du får hjälp av ett stort antal automatiska funktioner i %PRODUCTNAME Calc.  
Förutom de grundläggande räknesätten erbjuder %PRODUCTNAME Calc många beräkningsfunktioner som du kan mata in interaktivt med hjälp av Funktionsautopiloten.  
Med %PRODUCTNAME Calc kan du därför bekvämt utforma, fylla i, beräkna och skriva ut alla de formulär som du själv har skapat.  
Databasfunktioner  
Om dina data kan sammanfattas i dataposter, som t.ex. adresser, lagersaldon, kundorder eller dylikt, så kan du även förvalta dem med %PRODUCTNAME Calc.  
Även om du inte vill beräkna något, kan du t.ex. snabbt sortera databasområdet och söka efter vissa kännetecken i dina data som maximal - eller minimivärden.  
En tabell i %PRODUCTNAME Calc kan du dessutom använda som datakälla när du skapar standardbrev (kopplad utskrift) i %PRODUCTNAME Writer.  
Disponera data  
Du kan ordna data i översiktliga listor och visa dem i en viss ordning.  
Du behöver bara klicka några gånger med musen, så ordnas visningen så att t.ex. data i vissa områden visas eller döljs, formateras enligt speciella villkor eller del - och totalsummor beräknas.  
Undersöka data och göra prognoser  
Det finns många olika sätt att undersöka data som finns i %PRODUCTNAME Calc-tabeller. %PRODUCTNAME Calc är t.ex. ett effektivt hjälpmedel för alla som skriver ett examensarbete eftersom programmet även har flera statistiska funktioner som regressionsberäkning.  
Och även i vardagsarbetet har du hjälp av de inbyggda finansmatematiska funktioner na eftersom du t.ex. kan skriva ut utförliga tabeller för de löpande krediterna och lånen med dem.  
Vad-händer-om-beräkningar  
Särskilt intressant är möjligheten att ändra enstaka faktorer i en beräkning som är sammansatt av flera faktorer och sedan direkt se hur resultatet förändras av detta.  
Du kan t.ex. göra enkla ändringar av tidsperioden, räntesatsen eller avbetalningssummorna i en kreditberäkning och direkt se hur andra faktorer påverkas.  
Dessutom kan du förvalta mera omfattande tabeller i olika scenarion som utgår från sinsemellan olika villkor.  
Dynamiska diagram  
Med %PRODUCTNAME Calc är det lätt att strukturera data i tabellen på ett åskådligt sätt.  
Du markerar helt enkelt motsvarande data och klickar på ikonen Infoga diagram.  
Rita upp en ram på det önskade stället och gör inställningar för visningen av diagrammet i den dialogruta som öppnas.  
Diagrammet infogas på det valda stället och uppdateras dynamiskt när de data som diagrammet baserar på ändras.  
Dataimport och dataexport  
Du kan importera data från andra kalkylprogram, redigera dem i %PRODUCTNAME Calc och vid behov även exportera dem igen i andra exportformat.  
Datareferenser lokalt och i nätverket  
I stället för ett fast värde eller en matematisk formel som refererar till andra celler i tabellen, så kan varje cell i %PRODUCTNAME Calc även innehålla en referens till innehållet i andra dokument.  
De här dokumenten behöver inte ens ligga på hårddisken i din dator, de kan finnas på en annan dator i nätverket eller någonstans på Internet.  
Så hittar du den här funktionen...  
Menyn Redigera - Diagramdata  
Ikon på verktygslisten:  
Diagramdata  
Menyn Infoga - Rubrik...  
Menyn Infoga - Förklaring...  
Menyn Format - Förklaring... - fliken Placering  
Menyn Infoga - Dataetiketter...  
Menyn Format - Objektegenskaper... - Datapunkt / Dataserie - fliken Dataetiketter (vid dataserie och datapunkt)  
Menyn Infoga - Axlar...  
Menyn Infoga - Gitter...  
Ikoner på verktygslisten:  
Horisontellt gitter på / av  
Vertikalt gitter på / av  
Menyn Infoga - Statistik...  
Menyn Infoga - Specialtecken...  
Menyn Format - Objektegenskaper...  
Menyn Format - Objektegenskaper... - dialogrutan Datapunkt  
Menyn Format - Objektegenskaper... - dialogrutan Dataserie  
Menyn Format - Objektegenskaper... - dialogrutan Dataserie - fliken Alternativ  
Menyn Format - Rubrik  
Meny Format - Objektegenskaper... - dialogrutan Rubrik  
Menyn Format - Objektegenskaper... - dialogrutan Rubrik  
Menyn Format - Rubrik  
Menyn Format - Axel  
Menyn Format - Förklaring, Format - Objektegenskaper - dialogrutan FÃ¶rklaring  
Menyn Format - Axel  
Menyn Format - Axel - X-axel... eller Sekundär X-axel... eller Z-axel... eller Alla axlar...  
Menyn Format - Axel - Y-axel... eller SekundÃ¤r Y-axel...  
Menyn Format - Axel - Y-axel - fliken Skalning  
Menyn Format - Gitter  
Menyn Format - Gitter - X-, Y-, Z-axelhuvudgitter..., X-, Y-, Z-axelstÃ¶dgitter..., Alla axelgitter...  
Menyn Format - Diagramvägg - dialogrutan DiagramvÃ¤gg  
Menyn Format - Diagramgolv  
Menyn Format - DiagramomrÃ¥de  
Menyn Format - Diagramtyp  
Ikon på verktygslisten:  
Redigera diagramtyp  
Menyn Format - AutoFormat  
Ikon på verktygslisten:  
AutoFormat  
Menyn Format - 3D-vy  
Menyn Format - Placering  
Snabbmenyn Placering  
Rubrik på / av  
Axelrubrik på / av  
Horisontellt gitter på / av  
Axlar på / av  
Vertikalt gitter på / av  
Diagramdata  
Här öppnar du en dialogruta där du kan redigera diagrammets data.  
Dialogrutan är inte tillgänglig om du har infogat diagrammet i en %PRODUCTNAME Calc-tabell som visning av data i tabellen.  
Om du klickar på ikonen Diagramdata öppnas en dialogruta med många fler ikoner.  
Cellreferens  
I det här fältet visas cellreferensen i formen "kolumnbokstav + radnummer", t ex A1 för den första cellen i vänstra övre hörnet.  
Cellreferens  
Ignorera  
Det ersätts med det gamla innehållet.  
Ignorera  
Överta  
Klicka här om du vill överta inmatningsfältets ändrade innehåll i tabellen.  
Om du har gjort ett syntaxfel, så visas ett meddelande om detta.  
Då måste du korrigera felet i inmatningsfältet.  
Överta  
Inmatningsfält  
I inmatningsfältet visas det aktuella innehållet i den markerade cellen i tabellen och du kan redigera innehållet här.  
Tilldela  
Klicka på den här ikonen om du vill överföra tabellens data till diagrammet.  
Diagrammet uppdateras direkt med dessa nya data.  
Tilldela  
Infoga rad  
Klicka på den här ikonen om du vill infoga en ny tom rad ovanför den aktuella raden.  
Infoga rad  
Infoga kolumn  
Klicka här om du vill infoga en ny tom kolumn framför den aktuella kolumnen.  
Infoga kolumn  
Radera rad  
När Du klickar på den här ikonen, raderas den aktuella raden utan någon kontrollfråga.  
Den första raden med kolumnhuvudena kan Du inte radera.  
Radera rad  
Radera kolumn  
När Du klickar på den här ikonen, raderas den aktuella kolumnen utan någon kontrollfråga.  
Den första kolumnen med radrubrikerna kan Du inte radera.  
Radera kolumn  
Byt kolumner  
När Du klickar på den här ikonen, byts den aktuella kolumnens innehåll mot innehållet i kolumnen till höger om den.  
Ifall den sista kolumnen är utvald, så byts kolumninnehållet mot innehållet i den kolumn som står till vänster.  
Byt kolumner  
Byt rader  
Klicka på den här ikonen om Du vill byta den aktuella radens radinnehåll mot innehållet i den rad som ligger under den.  
Ifall den nedersta raden är utvald, så byts radinnehållet mot den näst sista radens radinnehåll.  
Byt rader  
Sortera kolumn  
Om Du vill att innehållet i den valda kolumnen ska sorteras stigande efter värde, så klickar Du på den här ikonen.  
Sortera kolumn  
Sortera rad  
Om Du vill att innehållet i den valda raden ska sorteras stigande efter värde, klickar Du på den här ikonen.  
Sortera rad  
Sortera tabellerna kolumnvis  
Klicka på den här ikonen om Du vill sortera tabellen kolumnvis.  
Hela datatabellen sorteras.  
Den aktuella kolumnen används som referens, sorteras och kolumnens övriga element flyttas i enlighet därmed.  
När sorteringen är klar, överförs databeståndet.  
Sortera tabellerna kolumnvis  
Sortera tabellerna radvis  
Klicka på den här ikonen om Du vill sortera tabellen radvis.  
Hela datatabellen sorteras.  
Den aktuella raden används som referens, sorteras och i enlighet därmed flyttas radens övriga element.  
När sorteringen är klar, överförs databeståndet.  
Sortera tabellerna radvis  
Diagramdatafält  
I huvudområdet i dialogrutan Diagramdata visas tabellen med data.  
Där finns rad - och kolumnhuvuden som hjälper dig att hitta rätt.  
Placera cellmarkören i den cell, rad eller kolumn som du vill redigera.  
I %PRODUCTNAME Chart kan du ångra flera redigeringssteg (antalet ställer du in under Verktyg - Alternativ - %PRODUCTNAME - Allmänt).  
Du kan visserligen även ångra redigeringen av diagramdata-tabellen stegvis, men resultatet visas i tabellen först när du har stängt dialogrutan Diagramdata en gång och öppnat den på nytt.  
Rubrik  
Här öppnar du en dialogruta där du kan skriva in och ändra texten i rubrikerna.  
Här väljer du hur huvudrubriken, underrubriken och rubrikerna för axlarna ska lyda och om de ska visas.  
Huvudrubrik  
Om Du aktiverar den här kryssrutan, kan Du skriva in den önskade huvudrubriken för objektet i textfältet.  
Underrubrik  
Om Du aktiverar den här kryssrutan, kan Du skriva in den önskade underrubriken i textfältet.  
Med ikonen Rubrik på / av på verktygslisten visar och döljer du huvud - och underrubriken.  
X-axel  
Om du aktiverar den här rutan, kan du skriva in den önskade rubriken för X-axeln i textfältet.  
Y-axel  
Om du aktiverar den här rutan, kan du skriva in den önskade rubriken för Y-axeln i textfältet.  
Z-axel  
Om du aktiverar den här rutan, kan du skriva in den önskade rubriken för Z-axeln i textfältet.  
Den här rutan kan du bara aktivera för tredimensionella diagram.  
Genom att klicka på ikonen Axelrubrik på / av på verktygslisten visar eller döljer du axelrubrikerna.  
Förklaring  
Här ändrar du placeringen av förklaringen i diagrammet.  
Med ikonen Förklaring på / av på verktygslisten kan du visa eller dölja förklaringen.  
Förklaring på / av  
Visa  
Aktivera den här rutan om du vill ha en förklaring till diagrammet. (Det här alternativet visas bara om du öppnar dialogrutan via Infoga - Förklaring.)  
Placering  
I det här området väljer du hur förklaringen ska visas.  
Till vänster  
Om du väljer det här alternativet, visas förklaringen till vänster om diagrammet.  
Uppe  
Om du väljer det här alternativet, visas förklaringen ovanför diagrammet.  
Till höger  
Om du väljer det här alternativet, visas förklaringen till höger om diagrammet.  
Nere  
Om du väljer det här alternativet, visas förklaringen nedanför diagrammet.  
Dataetikett  
Här öppnar du en dialogruta där du kan ställa in datapunkternas etiketter.  
Så kan du visa information om dina data.  
Dataetikett  
I det här området gör du dina val för dataetiketterna.  
Visa värde  
Klicka här om datapunkternas värden ska visas.  
I de tillhörande alternativfälten definierar du om värdet ska visas som tal eller i procent.  
som tal  
Markera den här rutan om du vill visa datapunkternas absoluta värden.  
i procent  
Markera det här alternativet om du vill visa den procentuella andelen för varje kolumns datapunkter.  
Visa etikettext  
Klicka här om du vill att beteckningen för datapunkterna ska visas.  
Visa förklaringssymbol bredvid etikett  
Klicka här om du vill placera symbolen som visas i förklaringen bredvid varje datapunktsetikett.  
Axlar  
Här bestämmer du vilka av axlarna som ska visas i diagrammet.  
Huvudaxel  
Markera den axel som ska visas i det här området.  
X-axel  
Markera den här rutan om X-axeln ska visas som linje med indelningsmärken.  
Y-axel  
Markera den här rutan om Y-axeln ska visas som linje med indelningsmärken.  
Z-axel  
Markera den här rutan om Z-axeln ska visas som linje med indelningsmärken.  
Den här axeln kan du bara visa i tredimensionella diagram.  
Sekundär axel  
I det här området kan du tilldela diagrammet en andra axel.  
Om en dataserie redan har tilldelats den här axeln, visar %PRODUCTNAME automatiskt axeln och etiketten.  
De här förinställningarna kan du stänga av i efterhand.  
Om det inte existerar någon tilldelning, och du aktiverar det här området, så övertas värdena för den primära axeln till den sekundära.  
X-axel  
Om du markerar den här rutan får diagrammet en andra X-axel.  
Y-axel  
Om du markerar den här rutan får diagrammet en andra Y-axel.  
Om du använder både huvudaxeln och den sekundära axeln kan du infoga skalning med olika finhet.  
Du kan till exempel skala en axel till 10 centimeter, den andra till 100 millimeter.  
Statistik  
Här bestämmer Du om Du vill visa statistikfunktioner, t ex medelvärde, felkategori eller regression, för 2D-objekt.  
Det här menykommandot kan Du bara välja för 2D-objekt.  
Medelvärde  
Om du markerar den här kryssrutan, visas det statistiska medelvärdet av dina diagramvärden.  
Felkategori  
I det här området kan Du välja bland de olika visningsformerna för respektive felkategori.  
Ingen funktion  
Välj detta alternativfält om Du inte vill ha någon visning.  
Varians  
Markera det här alternativfältet om Du vill visa en varians ur antalet datapunkter och de tillhörande värdena.  
Standardavvikelse  
Markera det här alternativfältet om Du vill visa en standardavvikelse (variansens kvadratrot).  
Procentuell  
Välj det här alternativfältet om Du vill ha en procentuell visning.  
Den här visningen gäller för respektive datapunkt.  
Ställ in det procentuella värdet i rotationsfältet.  
Största fel  
Markera det här alternativfältet om det största felet, med avseende på datagruppens största värde, ska visas i procent.  
Ställ in det procentuella värdet i rotationsfältet.  
Konstant värde  
Markera det här alternativfältet om Du vill visa det konstanta värdet i procent Ange det positiva värdet i rotationsfältet + och det negativa i rotationsfältet -.  
Felindikator  
I detta fält väljer du en felindikator.  
Du kan välja mellan Inga indikatorer, Indikatorer på båda sidor, Undre indikator och Övre indikator.  
Regressionskurvor  
Det här området är bara aktivt om Du har valt XY-diagram som diagramtyp.  
Välj mellan regressionskurvalternativen Ingen, Linjär, Logaritmisk, Exponentiell eller Potentiell regression.  
Alternativ  
I den här dialogrutan definierar du justering och avstånd för 2D-objekt.  
Justera dataserie mot:  
I det här området kan du välja mellan två skalningar av y-axeln.  
Axlarna kan bara skalas och förses med attribut separat.  
Primär Y-axel  
I standardinställningen är det här alternativet aktivt.  
Alla dataserier justeras efter den primära y-axeln.  
Sekundär Y-axel  
Om du vill ha en annan skalning av y-axeln, väljer du det här alternativfältet.  
Axeln syns bara om du tilldelar den minst en dataserie och visningen av axlarna inte är generellt avstängd.  
Inställningar  
Om du har skapat ett stapeldiagram med liggande staplar kan du göra inställningar i det här området.  
Alla ändringar gäller inte bara för den aktuella dataserien utan för alla dataserier i ditt diagram.  
Avstånd  
Här kan du ställa in avståndet mellan de enskilda kolumnerna med data i procent.  
Det största möjliga avståndet ligger på 600 Prozent.  
Överlappning  
Om dataserierna ska överlappa varandra kan du ställa in det i det här rotationsfältet.  
Du kan välja mellan -100 till +100 Prozent.  
Förbindelselinjer  
Vid stapeldiagram av typen "Staplat" och "Procent "förbinds nivåerna som hör ihop i alla kolumner med linjer om du klickar på den här rutan med musen.  
Gitter  
Du kan dela in axlarna med gitterlinjer.  
Som standard är bara y-axelns huvudgitter inkopplat.  
Huvudgitter  
I detta område fastställer Du för vilken axel Du vill ha ett huvudgitter.  
X-axel  
Markera det här fältet om Du vill att x-axeln ska grovindelas med gitterlinjer.  
Med ikonen Horisontellt gitter på / av på verktygslisten visar resp. döljer du gittret för x-axeln.  
Fältet Stödgitter får inte vara aktiverat.  
Stödgittret fortsätter alltså att visas.  
Y-axel  
Markera det här fältet om Du vill att y-axeln ska grovindelas med gitterlinjer.  
Med ikonen Vertikalt gitter på / av på verktygslisten visar eller döljer du gittret för y-axeln.  
Men förutsättningen är att fältet Stödgitter inte är aktiverat.  
Om du har aktiverat stödgittret kan du bara dölja huvudgittret.  
Stödgittret fortsätter att visas.  
Z-axel  
Markera det här fältet om Du vill att z-axeln ska grovindelas med gitterlinjer.  
Denna axel finns bara i 3D-diagram.  
Stödgitter  
Här kan Du infoga ett stödgitter för varje axel och därigenom ytterligare minska avstånden i indelningen.  
Det därtill hörande huvudgittret ska vara inkopplat.  
X-axel  
Markera det här fältet om Du vill att x-axeln ska finindelas med gitterlinjer.  
Y-axel  
Markera det här fältet om Du vill att y-axeln ska finindelas med gitterlinjer.  
Z-axel  
Markera det här fältet om Du vill att z-axeln ska finindelas med gitterlinjer.  
Denna axel kan bara infogas i 3D-diagram.  
Objektegenskaper  
Med det här kommandot tilldelar du det markerade objektet egenskaper.  
Beroende på vilket objekt du har markerat, öppnar du dialogrutor som du även når med följande kommandon på menyn Format:  
Diagramvägg...  
Diagramområde...  
Diagramgolv...  
Rubrik  
Förklaring...  
X-axel...  
Y-axel...  
Gitter  
Datapunkt  
Här ändrar du egenskaperna för en markerad datapunkt.  
Den här dialogrutan visas om du väljer menykommandot Format - Objektegenskaper när en enskild datapunkt är markerad.  
En del menykommandon är antingen bara tillgängliga till för 2D - eller 3D-diagram.  
Ändringarna som du gör här påverkar bara den aktuella datapunkten.  
Om du t.ex. ändrar färgen på en liggande stapel, så får bara den liggande stapeln en ny färg.  
Dataserie  
Här ändrar du egenskaperna för en markerad dataserie.  
Den här dialogrutan visas om du väljer menykommandot Format - Objektegenskaper när en dataserie är markerad.  
En del menykommandon är bara tillgängliga för 2D - eller 3D-diagram.  
Ändringarna som du gör här påverkar hela dataserien.  
Om du t.ex. ändrar färgen, så ändras alla element som hör till den här dataserien.  
Statistik  
Rubrik  
Det här menykommandot öppnar en undermeny där du kan ändra egenskaperna för rubrikerna i diagrammet.  
Huvudrubrik...  
Underrubrik...  
X-axelrubrik...  
Y-axelrubrik...  
Z-axelrubrik...  
Alla rubriker...  
Rubrik  
Här ändrar du egenskaperna för den markerade rubriken.  
Tecken  
Justering  
Under den här fliken kan du ändra justeringen av rubriketiketten.  
Det finns t.ex. skillnader mellan etiketteringen av 2D-objekt och 3D-objekt.  
Tänk på att det kan uppstå problem med att visa etiketteringen i diagram med för liten visningsstorlek.  
Du kan undvika detta genom att antingen förstora visningen eller minska teckenstorleken.  
Rubrik  
Här ändrar du egenskaperna för den markerade rubriken eller alla rubriker gemensamt.  
Tecken  
Etikett  
Under den här fliken kan du ändra justeringen av axeletiketten.  
Några av de listade alternativen är inte tillgängliga för alla etikettyper, det finns t.ex. skillnader mellan 2D - och 3D-objektetiketter.  
Visa etikett  
Om axeletiketterna inte ska visas, avmarkerar du den här rutan.  
Med den här ikonen på verktygslisten kan du visa och dölja etiketterna för alla axlar gemensamt.  
Rotera etikett  
I det här området kan du definiera skrivriktningen för cellinnehållet.  
För detta finns det två kommandoknappar som heter ABCD.  
ABCD  
Med hjälp av den runda kommandoknappen, som liknar en nummerskiva, kan Du steglöst och gradvis ställa in skrivriktningen med musen.  
Du får ett första synintryck genom att justeringen av tecknen ABCD ändrar sig efter Din inställning.  
ABCD  
Med den andra kommandoknappen kan Du bara ställa in en lodrät visning av cellinnehållet.  
En lodrät X-axeletikett kan komma att "klippas av" av X-axelns linje.  
Grader  
Under kommandoknapparna finns ett rotationsfält som du också kan använda för att definiera gradtalet.  
Textflöde  
I det här området kan Du bestämma textflödet för etiketterna.  
Överlappande  
Välj det här alternativet om axlarnas etiketter ska överlappa varandra.  
Detta kan vara lämpligt när det är ont om plats.  
För de olika titeljusteringarna finns inte detta alternativ.  
Brytning  
Markera den här kryssrutan om Du vill tillåta en brytning av texten.  
Följande alternativ är inte alltid tillgängliga:  
Placering  
Detta område kan Du bara välja om Du har skapat ett 2D-diagram och har öppnat menyn Format - Axel - Y-axel respektive X-axel.  
Här väljer Du hur axelns sifferetiketter ska placeras.  
Bredvid varandra  
Markera den här rutan om talen vid axeln vanligtvis ska placeras bredvid varandra.  
Upphöjt / nedsänkt  
Markera den här rutan om talen vid axeln ska placeras upphöjt och nedsänkt om vartannat.  
Nedsänkt / upphöjt  
Markera den här rutan om talen vid axeln ska placeras nedsänkt och upphöjt om vartannat.  
Automatiskt  
Markera den här rutan om talen vid axeln ska placeras automatiskt.  
Tänk på att det kan uppstå problem med visningen av etiketterna om diagrammet har för liten visningsstorlek.  
Du kan undvika detta genom att antingen förstora visningen eller minska teckenstorleken.  
Förklaring  
Här definierar du förklaringens inramning, yta, teckeneffekt och placering.  
Tecken  
Placering  
Axel  
Här öppnar du en undermeny där du kan ändra axlarnas egenskaper.  
Vilka flikar dialogrutorna innehåller beror på vilken diagramtyp du har valt.  
X-axel...  
Y-axel...  
Sekundär X-axel...  
Så snart Du har aktiverat denna extra X-axel under Infoga - Axlar, kan Du här bl a bestämma axelns linjestil, teckensnittet och skrivriktningen för axeletiketten.  
Sekundär Y-axel...  
Om Du tidigare har aktiverat denna extra Y-axel under Infoga - Axlar, kan Du här bl a bestämma axelns linjestil, teckensnittet och skrivriktningen för axeletiketten.  
Z-axel...  
Alla axlar...  
Axlar  
Med det här kommandot öppnar du en dialogruta där du kan ändra axel-egenskaperna.  
När du har valt alla axlar heter dialogrutan Axlar.  
För XY-diagram är även X-axelns dialogruta utökad med fliken Skalning.  
X-axeln kan bara skalas i diagramtypen XY.  
Tecken  
Y-axel  
Med det här kommandot öppnar du en dialogruta där du kan ändra axel-egenskaperna.  
När du har markerat alla axlar heter dialogrutan bara Axlar.  
Tecken  
Tal  
Skalning  
Under den här fliken styr du y-axelns skalning.  
I xy-diagram kan du även skala x-axeln här.  
Y-axeln skalas automatiskt av %PRODUCTNAME så att alla värden visas optimalt.  
Om du vill uppnå vissa effekter, kan du ändra axelskalningen för hand.  
Om du t.ex. inte visar staplarna i ett stapeldiagram i deras helhet, utan bara de övre delarna genom att flytta nollinjen uppåt, höjdskillnaderna mellan staplarna mer iögonfallande än om staplarna hade visats i sin helhet.  
Axelskalning  
I det här området anger du värdena för axelindelningen.  
De fem egenskaperna Minimum, Maximum, Huvudintervall, Hjälpintervall och Axel vid kan du låta sätta automatiskt.  
Minimum  
Ange ett nytt minimivärde för axelns startpunkt i det här textfältet.  
Maximum  
Ange ett nytt maximivärde för axelns slutpunkt i det här textfältet.  
Huvudintervall  
Här anger Du intervallet för axelns huvudindelning.  
Huvudintervallet får inte vara större än värdeområdet.  
Hjälpintervall  
Här anger Du intervallet för axelns hjälpindelning.  
Axel vid:  
Här anger Du den position utmed axeln där ursprunget för de visade värdena ska ligga.  
Om Du t ex har ett stapeldiagram där alla värden är större än noll, och lägger minimum på -10, så kan Du sedan även dra ned axeln till -10 och förlänga staplarna artificiellt på motsvarande sätt.  
Automatiskt  
Ta bort markeringen i en av rutorna Automatiskt, så kan du sedan ange ett nytt värde i textfältet.  
Om du vill arbeta med "fasta" värden bör du inaktivera det här alternativet.  
Detta förhindrar att det sker någon automatisk (dynamisk) skalning.  
Logaritmisk skalning  
Markera den här rutan om axeln ska indelas logaritmiskt.  
Använd denna funktion om du har värden som avviker kraftigt från varandra.  
Med logaritmisk skalning åstadkommer du att avstånden mellan axelns gitterlinjer är lika fastän de har olika värden.  
Axelmarkeringar  
I det här området kan du bestämma om markeringarna ska sättas på axelns in - eller utsida.  
Du kan även kombinera de båda alternativen.  
Detta leder till en heldragen markering som syns på insidan och på utsidan.  
inre  
Det här fältet anger att markeringen ligger på axelns insida.  
yttre  
Om du markerar det här fältet, så sätts markeringen på axelns utsida.  
Hjälpmarkeringar  
I det här området kan du definiera markeringsstreck mellan axelmarkeringarna.  
Detta innebär att en heldragen markeringslinje dras från utsidan till insidan.  
inre  
Aktivera det här fältet om hjälpmarkeringen ska ligga på axelns insida.  
yttre  
Aktivera det här fältet om hjälpmarkeringen ska ligga på axelns utsida.  
Gitter  
Detta kommando öppnar en undermeny där du kan välja vilket gitter som ska formateras.  
X-axelhuvudgitter...  
Y-axelhuvudgitter...  
Z-axelhuvudgitter...  
X-axelstödgitter...  
Y-axelstödgitter...  
Z-axelstödgitter...  
Alla axelgitter  
Gitter  
Här öppnar du dialogrutan Gitter där du definierar gitteregenskaperna.  
Diagramvägg  
Här ändrar du diagramväggens egenskaper.  
Diagramväggen är den "lodräta" bakgrunden bakom dataområdet i diagrammet.  
Diagramgolv  
Här ändrar du egenskaperna för diagramgolvet.  
Diagramgolvet är den undre ytan i tredimensionella diagram.  
Den här funktionen kan du därför bara välja för tredimensionella diagram.  
Diagramområde  
Här ändrar du egenskaperna för diagramområdet.  
Diagramområdet är bakgrunden bakom alla element i diagrammet.  
Diagramtyp  
Här kan du välja diagramtyp bland ett antal standardtyper.  
Diagramkategori  
Här anger Du om Du vill skapa ett tvådimensionellt eller tredimensionellt diagram.  
När Du har valt något av dessa alternativ, visas tillgängliga diagramtyper och tillhörande varianter.  
2D  
Om Du markerar det här alternativet, kan Du sedan välja bland de tvådimensionella diagramtyperna i fälten Typ och Variant.  
3D  
Om Du markerar det här alternativet, kan Du sedan välja bland de tredimensionella diagramtyperna i fälten Typ och Variant.  
Du kan välja ytterligare alternativ via 3D-effekter på menyn Format.  
Du kan även rotera 3D-diagram interaktivt.  
Om Du klickar på diagrammet visas en böjd markörpil vid vilken objektet kan roteras runt sina axlar.  
Diagramtyp  
Här kan du välja mellan alla tillgängliga diagramtyper.  
Urvalet omfattar alla vanliga typer inklusive XY-diagram och polärdiagram.  
Den markerade typen visas inramad och namnet visas i den nedre delen av området.  
I kategorin 2D-diagram har du tillgång till linjer, ytor, staplar, liggande staplar, cirklar, XY-diagram, polär - och kursdiagram.  
Polär-, XY - och linjediagram visas med grå bakgrund, vilket förbättrar visningen rent optiskt.  
Den här standardinställningen kan du givetvis ändra.  
I de s.k. tårtdiagrammen (cirkeldiagram i form av en tårta) kan du dra ut de enskilda tårtbitarna med musen.  
Då ändras radien för alla bitar eftersom hela diagrammet visas i en ram med förinställd storlek.  
Men du kan markera diagrammet sedan och ändra dess storlek.  
I kursdiagram används symboler för att markera kursernas rörelse uppåt och nedåt, omsättningar och det totala antalet aktier.  
Dessa symboler har som standard en storlek som inte överstiger linjebredden.  
På så vis blir punkterna så att säga osynliga.  
Endast slutkursen markeras med ett synligt streck.  
Först om Du själv integrerar andra grafiska objekt blir alla punkter synliga.  
I kategorin 3D-diagram kan du välja typerna linjer, ytor, staplar, liggande staplar och cirklar.  
Om du vill välja en viss typ behöver du bara klicka på bilden.  
Samtidigt visas de tillhörande varianterna i området Variant.  
Om Du ändrar axelgraderingen för linje-, yt - och XY-diagram, och några symboler ligger utanför gittret, så kan detta medföra att visningen blir ofullständig.  
Även statistiklinjer visas bara om deras centrum ligger inom rektangelområdet.  
Variant  
Här visas diagramtypernas varianter, och du kan välja en av dem.  
De tillgängliga varianterna skiljer sig åt beroende på vilken dimension och diagramtyp du väljer.  
Om du t.ex. har valt 2D-stapeldiagrammet kan du använda varianterna Normal, Staplat, Procent och Kombinationsdiagram.  
Om du vill visa ditt diagram som liggande 3D-staplar, kan du bl.a. välja bland olika rör - pyramid - och konvarianter.  
Den variant som du väljer gäller för hela diagrammet.  
Om Du har aktiverat kommandot Tips på menyn Hjälp och sedan placerar muspekaren ovanför ikonerna, så visas namnen både för diagramtyperna och för deras varianter.  
Även om Tips-hjälpen inte är aktiverad, så visas åtminstone namnet för den markerade typen respektive den markerade varianten i det tillhörande området.  
Punktordning  
Vid linjediagram och XY-diagram kan Du välja en av spline-varianterna.  
Du ser det här rotationsfältet vid B-splines.  
Här bestämmer Du ordningen för B-splinekurvan.  
Vid 1 är resultatet en linje, vid 2 en parabel, vid n i allmänhet en parabel av n-ordning.  
Upplösning  
Vid linjediagram och XY-diagram kan Du välja en av spline-varianterna.  
Då visas det här rotationsfältet.  
Här bestämmer Du antalet beräknade mellanpunkter på spline-kurvan mellan två datapunkter.  
AutoFormat  
Med det här kommandot öppnar du dialogrutan AutoFormat diagram.  
På sidorna i dialogrutan kan du ändra många av diagrammets egenskaper interaktivt.  
<< Tillbaka  
I dialogrutan kan Du titta på förhandsvisningen av det föregående arbetssteget.  
Aktuella inställningar bibehålls.  
Denna kommandoknapp är endast tillgänglig fr o m andra redigeringssteget.  
Nästa >>  
Om du klickar på den här kommandoknappen använder %PRODUCTNAME de aktuella inställningarna i dialogrutan och går vidare till nästa redigeringssteg.  
Om du har kommit till den sista sidan i dialogrutan går det inte att klicka på den här kommandoknappen.  
Färdigställ  
%PRODUCTNAME skapar ett nytt diagram baserat på dina inställningar.  
3D-vy  
Här anger Du perspektivvinkeln för 3D-diagrammet i det tredimensionella rummet.  
Det här menykommandot är bara tillgängligt om Du har valt ett 3D-diagram som diagramtyp.  
Axelrotation  
Här anger Du vinklarna för axelrotationen.  
X-axel  
Här anger du rotationsvinkeln runt X-axeln från vilken du vill titta på diagrammet.  
Med vinkeln 0 grader tittar du på diagrammet direkt från X-axelns höjd, med vinkeln 90 grader direkt uppifrån.  
Y-axel  
Här anger du rotationsvinkeln runt Y-axeln från vilken du vill titta på diagrammet.  
Med vinkeln 0 grader tittar du på diagrammet direkt framifrån, med vinkeln 90 grader direkt från höger sida.  
Z-axel  
Här anger du rotationsvinkeln runt Z-axeln från vilken du vill titta på diagrammet.  
Med vinkeln 0 grader tittar du på diagrammet i normalläge, med vinkeln 90 grader tippar du diagrammet så att säga på den vänstra sidan.  
Axelrotationen runt Z-axeln är inte tillgänglig för alla tredimensionella diagram.  
Placering  
Här kan du ändra ordningsföljden för diagrammets dataserier i efterhand.  
Dataposternas positioner i datatabellen förblir oförändrade.  
Du kan bara använda kommandona när du infogar ett diagram i %PRODUCTNAME Calc.  
Den här funktionen kan du bara använda om du visar data kolumnvis.  
Du kan inte byta till radvis visning.  
Längre fram  
På detta sätt flyttar Du den markerade dataserien i diagrammet längre fram (åt höger).  
Längre bak  
Med det här kommandot förskjuter Du den markerade dataserien i diagrammet bakåt (åt vänster).  
Data i rader  
Här ändras tilldelningen av data för diagrammet.  
Det innebär att först visas de data bredvid varandra som står i kolumn 1, till höger om dem visas sedan de data som står i kolumn 2 o.s.v.  
Data i rader  
Data i kolumner  
Här ändras tilldelningen av data för diagrammet.  
Det innebär att först visas de data bredvid varandra som står på rad 1, till höger om dem visas sedan de data som står på rad 2 o.s.v.  
Data i kolumner  
Textskalning  
Här aktiverar du textskalningen.  
Om du har aktiverat textskalningen (ikonen är intryckt) och ändrar storleken på fönstret där diagramobjektet finns, så ändras samtidigt texternas storlek.  
Om textskalningen inte är aktiverad, behåller texterna sin storlek.  
Textskalning  
Ordna diagrammet på nytt  
Om du klickar på den här ikonen återställs den ursprungliga visningen av diagrammet.  
Ordna diagrammet på nytt  
Aktuell diagramtyp  
I det här fältet på statuslisten visas den aktuella diagramtypens namn.  
Diagram i %PRODUCTNAME  
I %PRODUCTNAME kan du infoga diagram i dina dokument.  
Information om diagramfunktioner  
Referenshjälp  
Menyerna för diagram  
Symbollisterna för diagram  
Menyer  
När du arbetar med diagram hittar du kommandon för att öppna de olika programfunktionerna på menylisten.  
Kommandon på snabbmenyn  
Redigera  
Växlar till redigeringsläge.  
Arkiv  
På den här menyn hittar du kommandon som används till att hantera och skriva ut dokument och avsluta tillämpningen.  
Öppna...  
Spara som...  
Versioner...  
Dokument som e-post...  
Egenskaper...  
Skriv ut...  
Skrivarinställning...  
Redigera  
Här hittar du diagramdata för det markerade diagrammet.  
Visa  
På den här menyn kan du bland annat visa och dölja symbollister och statuslisten.  
Infoga  
Här finns kommandon som används till att infoga rubriker, förklaringar, dataetiketter, axlar och gitter samt statistikfunktioner.  
Rubrik...  
Förklaring...  
Dataetiketter...  
Axlar...  
Gitter...  
Statistik...  
Specialtecken...  
Bara tecken som finns i det aktuella teckensnittet är tillgängliga.  
Format  
På den här menyn definierar du utseendet för diagramdokument.  
Du kan styra alla aspekter av diagrammets utseende i olika dialogrutor och på olika undermenyer.  
Objektegenskaper...  
Förklaring...  
Diagramvägg...  
Diagramgolv...  
Diagramområde...  
Diagramtyp...  
AutoFormat...  
3D-vy...  
Verktyg  
På den här menyn hittar du kommandon som används till att anpassa gränssnittet och göra standardinställningar för programmet.  
Anpassa...  
Fönster  
På fönstermenyn kan du öppna fönster.  
Där finns även en lista över öppna dokument.  
Symbollister  
Här finns beskrivningar av ikonerna på verktygslisten, som används till att utföra de vanligaste kommandona.  
Statuslist  
På statuslisten visas aktuell information om dokumentets status.  
Verktygslist  
Verktygslisten är placerad i vänstra kanten av diagramfönstret.  
Där har du tillgång till viktiga funktioner som du ofta behöver.  
Rubrik  
Förklaring  
Axelrubrik  
Axlar  
Horisontellt gitter  
Vertikalt gitter  
Överblick över %PRODUCTNAME Chart  
Här ger vi dig en kort överblick över de omfattande diagramfunktionerna i %PRODUCTNAME.  
I ett tabelldokument eller i en tabell i ett textdokument kan du markera ett område med data och sedan infoga ett diagram direkt med dessa data.  
Data i det markerade området överförs till diagrammet med en "levande" förbindelse.  
Det betyder att diagrammet ändras automatiskt när de data som används för diagrammet ändras i dokumentet.  
Många diagramtyper  
Välj bland normala tvådimensionella diagram, t.ex. stapeldiagram, kurvdiagram, kursdiagram, eller välj 3D-diagram, där du kan använda många möjligheter till optisk anpassning.  
Du kan lätt byta från en diagramtyp till en annan.  
När det gäller kurvdiagram kan du visa många statistiska egenskaper, som %PRODUCTNAME beräknar.  
Det finns fyra varianter av kursdiagram.  
Du kan bland annat skapa kombinationer av omsättning och typiska kursdata.  
I %PRODUCTNAME kan du visa ett valfritt antal dataserier som kursdiagram.  
För många diagramtyper kan du infoga hjälpmarkeringar intill de egentliga markeringarna på axellinjerna för att uppnå bättre skalning.  
Universella formateringar  
Du kan formatera de enskilda elementen i diagrammen via snabbmenyerna respektive de normala menyerna och symbollisterna.  
Du kan bl.a. göra långtgående anpassningar av bildtext, skalning, bakgrund och andra element efter dina önskemål om hur ett diagram ska se ut.  
Så hittar du den här funktionen...  
Sida  
Om du väljer det här kommandot infogas en ny tom sida i dokumentet.  
Om det finns fler sidor flyttas de bakåt och får nya standardnamn.  
Om du t.ex. infogar en sida efter Sida 2 så kommer Sida 3, om den finns, att heta Sida 4.  
Kortkommandon för teckningsdokument  
Här hittar du en lista med tangentkombinationer som du kan använda i teckningsdokument.  
Dessutom gäller de allmänna tangentkombinationerna i %PRODUCTNAME.  
Funktionstangenter vid teckningsdokument  
Tangentkombination  
Effekt  
F2  
Redigera text  
F3  
Gå in i gruppering  
Kommando Ctrl +F3  
Lämna gruppering  
Skift+F3  
Dialogrutan Duplicera  
F4  
Dialogrutan Position och storlek  
F5  
Navigator  
F7  
Rättstavningskontroll  
Kommando Ctrl +F7  
Synonymordlista  
F8  
Redigera punkter på / av  
Kommando Ctrl +Skift+F8  
Anpassa text till ram  
F11  
Stylist  
Tangentstyrning i teckningsdokument  
Tangentkombination  
Effekt  
+ tangent  
Förstorar vyn  
- tangent  
Förminskar vyn  
×-tangent (numeriska delen av tangentbordet)  
Zoom på hela sidan  
÷-tangent (numeriska delen av tangentbordet)  
Zoom till den aktuella markeringen  
Skift + Kommando Ctrl +G  
Gruppering  
Skift + Kommando+Alternativ Ctrl+Alt +A  
Upphäv gruppering  
Skift + Kommando Ctrl +K  
Kombination  
Skift + Kommando+Alternativ Ctrl+Alt +K  
Upphäv kombination  
Skift + Kommando Ctrl +( plustecken)  
Längst fram  
Kommando Ctrl +( plustecken)  
Längre fram  
Kommando Ctrl -( minustecken)  
Längre bak  
Skift + Kommando Ctrl -( minustecken)  
Längst bak  
Speciella tangentstyrningar vid teckningsdokument  
Tangentkombination  
Effekt  
Piltangent  
Flyttar det markerade objektet i pilens riktning  
Kommando Ctrl +piltangent  
Flyttar sidvyn i önskad riktning.  
Nedtryckt skifttangent och dra med musen  
Det markerade objektet flyttas exakt horisontellt eller vertikalt i den önskade riktningen.  
Kommando Ctrl och dra med musen med alternativet Kopia vid förflyttning aktivt  
När du flyttar det markerade objektet skapas en kopia.  
Alternativ Alt  
När du skapar eller ändrar storlek på objekt, centreras de om du först trycker på tangenten Alternativ Alt.  
Alternativ Alt och klicka med musen på objekt  
Markering av objekt som överlappar varandra.  
Objektet som ligger bakom det markerade objektet markeras.  
Alternativ Alt +Skift och klicka med musen på objekt  
Markering av objekt som överlappar varandra.  
Objektet som ligger framför det markerade objektet markeras.  
Skifttangent vid markering  
Objekt läggs till markeringen om det ännu inte markerats eller tas bort från markeringen om det redan varit markerat innan.  
Skifttangent vid förstora / skapa  
Objektet förstoras proportionellt mot ursprungsformen.  
En rak linje kan bara ändras i sin riktning.  
Tabbtangent  
De enskilda objekten markeras i den ordning de skapades, från det första till det sista objektet.  
Skift+tabbtangent  
Markering av objekten i den ordning de skapades, från det sista till det första objektet.  
Skifttangent när du drar med musen i läget Redigera punkter  
Gör det möjligt att ändra längden på en måttlinje.  
Esc-tangent  
Skiftar till markeringsläget när ett skapa-verktyg är aktivt.  
Avmarkerar ett markerat objekt.  
Stänger av textinmatningsläget för ett objekt som står i textinmatningsläget.  
Objektet fortsätter att vara markerat  
Placera och justera objekt  
Placering av objekt  
Om dina objekt överlappar varandra och du vill sätta enstaka objekt i förgrunden eller i bakgrunden, kan du antingen använda snabbmenyn eller ikonerna på utrullningslisten Placering.  
Klicka på ett objekt vars position du vill ändra i placeringen framför / bakom andra objekt.  
Klicka sedan på en av ikonerna i den övre raden på utrullningslisten Placering för att t.ex. placera objektet längst bak.  
Om du vill placera det bakom ett objekt, kan du klicka på ikonen Bakom objektet.  
Sedan klickar du på objektet bakom vilket det aktuella objektet skall placeras.  
En effekt ser du naturligtvis bara om objekten överlappar varandra nu eller när du har flyttat dem.  
Då byter objekten plats med varandra.  
Justering av objekt  
Objekten kan du dra med musen till varje position.  
Om du vill placera ett objekt precis vid övre sidmarginalen eller två objekt exakt vertikalt centrerade ovanför varandra, är det enklare att använda ikonerna på utrullningslisten Justering.  
Markera ett enskilt objekt och klicka sedan på en av ikonerna på utrullningslisten Justering.  
Objektet justeras då vid sidmarginalerna.  
Om du har markerat två eller fler objekt samtidigt justeras de till varandra.  
En särskild typ av justering är fördelning av objekt.  
Om du markerar minst tre objekt samtidigt, kan du använda kommandot Fördelning.  
I %PRODUCTNAME Impress och %PRODUCTNAME Draw hittar du kommandot på snabbmenyn, i %PRODUCTNAME Draw även på menyn Ändra.  
De markerade objekten fördelas så att deras kanter eller mittpunkter har samma avstånd från varandra.  
De båda objekten som är längst från varandra horisontalt resp. vertikalt, gäller som ej flyttbara fixpunkter.  
De andra objekten mellan de yttre objekten kan flyttas med den här funktionen.  
Tänk på att du har en ångra-funktion i flera nivåer överallt i %PRODUCTNAME.  
Aktivera den här funktionen genom att till exempel klicka på ikonen Ångra på funktionslisten eller genom att trycka på Kommando Ctrl +Z.  
För varje gång du väljer kommandot ångrar du en funktion.  
Definiera egna färger  
Du kan definiera ett valfritt antal egna färger, namnge dem och arkivera dem i färgpalettfiler.  
Välj Format - Yta i ett teckningsdokument.  
Dialogrutan Yta öppnas.  
Klicka på fliken Färger i dialogrutan.  
Här hittar du allt som du behöver för att ändra färgen på det aktuella objektet, men du kan också definiera och administrera fler färger här.  
Om du vill ge det aktuella dokumentet en ny färg som inte finns med i färgtabellen ännu, måste du först definiera den här nya färgen och ge den ett eget namn.  
De sparas automatiskt och går inte att ångra.  
Det kan däremot uppstå problem om du ändrar standardfärgerna.  
När en ny färg skall definieras är det bäst att först välja ut en färg som liknar den nya färgen i färgtabellen.  
Den visas för jämförelse i det övre förhandsvisningsfältet.  
I listrutan väljer du sedan färgmodell enligt vilken du vill definiera den nya färgen.  
I listrutan finns alternativen RGB och CMYK.  
Färgmodellerna RGB och CMYK hör till de mest använda modellerna för att definiera färger.  
RGB står för Rött-Grönt-Blått och beskriver de motsvarande färgandelarna, om färgerna på datorskärmen sammansätts utifrån de tre grundfärgerna.  
CMYK står för Cyan-Magenta-Yellow-blacK eller Cyan-Magenta-Yellow-Key och är färgmodellen som beskriver den subtraktiva färgproduktionen med utskriftsfärger.  
Välj färgmodellen som motsvarar det önskade utmatningsmediet (bildskärm eller skrivare).  
Om du lämnar bildfiler för fotografering är det bäst att fråga kopieringsservicen vilken färgmodell och vilket format de använder.  
Ställ in färgen genom att ändra värdena i rotationsfälten.  
Du kan mata in värden eller klicka på pilknapparna för att ändra de visade värdena.  
I det undre förhandsvisningsfältet ser du genast effekten.  
Du ser då dialogrutan Färg.  
Välj färg och stäng dialogrutan med OK.  
Om du tycker om färgen måste du nu bestämma om den nya färgen skall ersätta ursprungsfärgen eller om den skall definieras oberoende av ursprungsvärdet.  
Klicka på Ändra om du vill ersätta den bestående färgen som visas i det övre förhandsvisningsfältet.  
Du bör bara göra detta med färger som du har definierat själv.  
För att definiera den nya färgen matar du först in ett nytt namn i fältet Namn, klickar sedan på Lägg till och OK.  
Din nya färg är genast tillgänglig tillsammans med de andra färgerna.  
Om du stänger dialogrutan med Avbryt färgas inte det aktuella objektet om, men ändringarna av färgtabellen gäller i alla fall.  
Det finns mer information om att spara och ladda färgpaletter och andra palettfiler i %PRODUCTNAME -hjälpen.  
Färglist  
Kombinera objekt och bilda former  
I %PRODUCTNAME Draw och %PRODUCTNAME Impress kan du kombinera grafiska objekt på olika sätt.  
Det går att skapa nya objekt av flera enskilda objekt genom att använda logiska mängdoperatorer på ursprungsgeometrin.  
Kombinera objekt  
Markera flera objekt.  
Välj Kombinera på snabbmenyn.  
I motsats till gruppering där bara enskilda objekt sammanfogas, sammanfogar en kombination delobjekt till ett enda nytt geometriskt objekt med nya egenskaper.  
Kombinationen kan upphävas igen senare, men delobjektens enskilda attribut går förlorade.  
Den mest iögonfallande egenskapen hos en kombination ser du när de enskilda objekten överlappar varandra.  
I det här fallet stansas snittmängden ut som "hål" på alla ställen där ett antal objekt överlappar varandra.  
Detta är ett logiskt exklusiv-ELLER (XOR).  
På bilden ser du några objekt innan de kombineras till vänster, efter att de har kombinerats till höger.  
Kombinationens attribut hämtas från det objekt som står längst bak.  
Bilda former  
Kommandona Former - Sammansmält, Dra ifrån och Skär av bildar också ett nytt geometriskt objekt av de ursprungliga objekten.  
Det nya objektet uppstår genom att logiska mängdoperatorer används på den ursprungliga geometrin.  
Markera flera objekt.  
Välj Former på snabbmenyn.  
På undermenyn väljer du Sammansmält, Dra ifrån eller Skär av.  
På de följande bilderna ser du de ursprungliga ytorna till vänster och resultatet av kommandot bredvid till höger.  
Former - Sammansmält  
De markerade polygonerna smälts samman så att du får ett objekt vars yta är summan av alla delobjekt (logiskt ELLER).  
Former - Dra ifrån  
Alla andra markerade polygoner dras ifrån den polygon som ligger underst.  
Då bildas en sammansmältning av de andra polygonerna, sedan dras den ifrån polygonen som är placerad längst bak.  
Det tas hänsyn till hål.  
Logiskt motsvarar den här operationen följande formel:  
A - (B1 _BAR_..... _BAR_ Bn)  
Former - Skär av  
De markerade polygonerna sammanfattas till en enda polygon som motsvarar snittmängden av alla ytor (logiskt OCH).  
Bara de ytor blir över där alla polygoner överlappar varandra.  
Använd t.ex. även Former - Dra ifrån och Former - Skär av om du ska skära ut delar av en bitmapgrafik.  
Bilden innehåller exempel.  
Tona över mellan två objekt  
Det går bara att tona två objekt i teckningsdokument i %PRODUCTNAME Draw och inte i %PRODUCTNAME Impress.  
Om du behöver ett objekt med en toning i en presentation kan du kopiera det från teckningsdokumentet till presentationsdokumentet via urklippet.  
Vid toning beräknas en övergång mellan två objekt och övergångsnivåerna placeras på sidan.  
I övergångsnivåerna anpassas bland annat formen, orienteringen och färgen på objekten jämnt till varandra.  
Rita till exempel ett objekt nere till vänster i ett tomt teckningsdokument och ett annat objekt uppe till höger (välj olika färger).  
Markera båda objekten.  
Du kan nu göra fler inställningar i en dialogruta.  
Klicka på OK.  
%PRODUCTNAME Draw beräknar nu övergångsnivåerna och visar dem.  
Det här nya objektet är en gruppering som består av det ovannämnda antalet enskilda objekt.  
Du kan gå in i grupperingen (F3) och sedan redigera de enskilda objekten.  
Kommandona för arbete med grupperingar hittar du på menyn Ändra i %PRODUCTNAME Draw, under Format - Grupp eller på snabbmenyn i %PRODUCTNAME Impress.  
Det finns mer information i %PRODUCTNAME -hjälpen.  
Redigera - Tona över  
Rita sektorer och segment  
På utrullningslisten Ellipser ser du också ett antal ikoner som du kan använda om du vill rita sektorer och segment.  
Sektorer ser ut som perfekta "tårtbitar".  
Segment liknar bitarna som man får om man delar en tårta på mitten.  
Att teckna en ellips - eller cirkelsektor är en process i flera steg:  
1.  
Öppna utrullningslisten Ellipser och klicka på ikonen Cirkelsektor, ofylld.  
Markören blir ett hårkors med en liten sektor.  
2.  
Dra med nertryckt musknapp.  
Konturen av en cirkel följer musens rörelser.  
Första gången du klickar definierar du det första hörnet i en begränsningsrektangel som omsluter den ritade cirkeln.  
Begränsningsrektangeln känner du igen senare när du markerar cirkeln på de åtta handtagen i hörnen och på sidornas mitt.  
Om du hellre vill rita cirkeln från mitten så att det första klicket definierar dess mitt, så håller du ner Alternativ Alt -tangenten medan du drar.  
3.  
Släpp musknappen när cirkeln är så stor som du vill ha den.  
Nu ser du att en radie ritas i cirkeln som följer varje musrörelse.  
4.  
Placera radien så som den ena kanten av sektorn skall ligga och klicka sedan en gång.  
5.  
När du nu rör musen är den första radien definierad och en andra radie följer musens rörelse.  
Så fort du klickar igen är cirkelsektorn färdig.  
Du gör likadant när du ritar ellipssektorer.  
Genom måtten på begränsningsrektangeln som du drar upp i steg 2, bestämmer du ellipsens mått.  
Om du ritar ett segment gör du på samma sätt som beskrevs ovan för sektorerna.  
Det är inte en andra radie som följer musens rörelse utan en sekant genom cirkeln.  
Det finns fler ikoner på utrullningslisten Ellipser som du kan rita ellips - och cirkelbågar med.  
Även detta sker på samma sätt som beskrivs ovan, men i det här fallet ritas bara ellipsens eller cirkelns omfång.  
Duplicera objekt  
Duplicering av objekt gör det möjligt att enkelt skapa ett definierat antal kopior av ett objekt, som skiljer sig åt i position, orientering, storlek och färg från en kopia till en annan.  
Om du till exempel behöver en stapel med mynt kan du dra nytta av dupliceringsfunktionen.  
Det enda du behöver göra är att skapa det understa myntet:  
1.  
Rita en ellips eller en cirkel vid den undre sidmarginalen.  
2.  
Välj Redigera - Duplicera.  
Du ser dialogrutan Duplicera.  
3.  
Mata in följande värden:  
4.  
Välj ungefär 30 som antal kopior.  
X-axeln är den horisontala axeln från vänster till höger; förskjutning med positiva värden har en förskjutning åt höger till följd.  
Om myntstapeln skall växa nerifrån och upp, så måste du ange en negativ förskjutning i Y-riktningen.  
5.  
Om mynten skall bli mindre längre upp så matar du in ett negativt tal för bredd och höjd som förstoringsvärde.  
6.  
Nu återstår bara att mata in ändringen av färgerna nerifrån och upp.  
Välj till exempel en något mörkare gul som startfärg än för slutfärgen.  
7.  
Klicka på OK så skapas kopiorna.  
Redigera - Duplicera  
Ersätta färger med pipetten  
Du kan redigera infogade bilder i ett bitmapformat (t.ex. GIF, JPG) och metafilbilder (t.ex. WMF) med pipett en i %PRODUCTNAME Draw och %PRODUCTNAME Impress.  
Aktivera pipetten med kommandot Verktyg - Pipett.  
Du ser sedan fönstret Pipett.  
Pipetten kan ersätta utvalda färger och liknande färger i ett toleransområde med andra färger.  
Du kan ersätta upp till fyra färger samtidigt.  
Om du inte tycker om ersättningen kan du återställa allt genom att klicka på Ångra på funktionslisten.  
Använd pipetten för att t.ex. anpassa färgerna på olika bitmaps till varandra eller för att ge en bitmap färgerna från din företagslogotyp.  
Även attributet Transparens gäller som färg.  
Du kan ersätta transparensen i en bild med en färg, t.ex. med vitt.  
Det kan vara till hjälp om t.ex. din skrivardrivrutin har problem med att skriva ut transparenta grafikobjekt.  
Om du producerar en bild för publicering på HTML-sidor på Internet, t.ex. en bild på en produkt, gör det ofta ett bättre intryck om bilden inte är fyrkantig, utan bara innehållet är synligt mot webbsidans bakgrund.  
Om produkten har en vit bakgrund på bilden använder du pipetten för att ersätta färgen vitt med transparent och sparar resp. exporterar bilden i ett format som tillåter transparens (som t.ex. GIF).  
Vid den här metoden bör produkten naturligtvis inte ha några vita delar eftersom de skulle bli lika genomskinliga som bildens bakgrund.  
Så ersätter du färger med pipetten  
Infoga en bild i ett bitmap-format (t.ex. BMP, GIF, JPG, TIF) eller i ett metafilformat (t.ex. WMF).  
Välj Infoga - Grafik i %PRODUCTNAME Draw och %PRODUCTNAME Impress.  
Öppna fönstret Pipett via kommandot Verktyg - Pipett.  
Klicka på pipettikonen uppe till vänster i fönstret Pipett.  
Muspekaren blir till en särskild pekare som du kan använda till att peka på färgen som skall ersättas i det aktuella dokumentet.  
Färgfältet i fönstret Pipett visar färgen som är under muspekaren.  
Klicka med den vänstra musknappen när du har hittat färgen som skall ersättas.  
Den här färgen förs automatiskt in i den första av de fyra raderna i fönstret Pipett.  
I listrutan till höger på samma rad väljer du ut den nya färgen som skall ersätta den markerade färgen i hela bitmapbilden.  
Om du vill ersätta en färg till i samma bearbetningssteg, kan du klicka på rutan framför nästa rad, sedan på pipettikonen uppe till vänster igen och välja en färg på nytt.  
Det är möjligt att redigera upp till fyra färger samtidigt.  
Klicka på bitmapbilden eller metafilbilden där du vill ersätta färgerna så att den är markerad.  
Klicka på Ersätt i fönstret Pipett.  
Om för många liknande färger har ersatts kan du ångra steget, t.ex. med Kommando Ctrl +Z och minska färgtoleransen i rotationsfältet.  
Sedan klickar du på Ersätt igen.  
Pipett  
Definiera färggradient  
Om du vill tilldela ett objekt en färggradient från urvalet av redan definierade färggradienter, gör du så här:  
Markera objektet.  
Välj Yta på snabbmenyn eller på menyn Format.  
Välj alternativet Färggradient och sedan väljer du från listan över färggradienter.  
Så här definierar du en egen färggradient  
Du kan definiera en egen färggradient, spara den aktuella färggradienttabellen som fil eller ladda en annan tabell från en fil.  
Om du har markerat ett objekt och sedan definierar en ny gradient, tilldelas den nya gradienten genast det markerade objektet.  
Om du inte vill detta måste du upphäva markeringen innan du öppnar dialogrutan där färggradienter definieras.  
Klicka med urvalsverktyget på ett ställe där det inte finns något objekt.  
1.  
Klicka på fliken Färggradienter i dialogrutan Yta.  
Här väljer du alternativ för nya gradienter.  
2.  
Välj en gradient som du vill använda som utgångspunkt för din nya gradient i listan med gradienter och klicka på den.  
3.  
Klicka på Lägg till.  
Du ser en dialogruta där du kan mata in ett namn för den nya gradienten.  
I exemplet har vi matat in "Ufo" och klickat på OK.  
I slutet av listan finns det nu en ny post med det nya namnet som redan är markerad för redigering.  
4.  
Klicka på Ändra för att spara ändringarna i den nya gradienten.  
I förhandsvisningsfältet ser du hur gradienten kommer att se ut.  
5.  
Stäng dialogrutan med OK.  
Du kan börja använda den nya färggradienten direkt.  
Så här ändrar du en färggradient interaktivt  
Du kan ändra färggradienter genom att klicka och dra med musen.  
Förutsättning för att kunna definiera en färggradient interaktivt är att objektet redan har en färggradient.  
1.  
Markera ett objekt som innehåller en färggradient.  
2.  
Öppna utrullningslisten Effekter på verktygslisten i %PRODUCTNAME Draw.  
3.  
Klicka på ikonen Färggradient på utrullningslisten Effekter.  
Du ser nu två färgobjekt som är ihopkopplade med en vektor.  
Beroende på typ av färggradient kan du flytta ett eller båda färgobjekten med musen och definiera ursprung, slut och vinkel för färggradienten.  
Om du har öppnat färglisten, kan du dra färger till varje färgobjekt per dra-och-släpp för att på så sätt definiera start - och slutfärg.  
På samma sätt kan du definiera transparensen för ett objekt med hjälp av ikonen Transparens.  
Här definierar du en gråskalegradient från svart (0% transparens, täckande) till vitt (100% transparens, genomskinlig).  
Infoga grafik  
Välj kommandot Infoga - Grafik.  
Dialogrutan Infoga grafik öppnas.  
Välj grafikobjekt och klicka på Öppna.  
Markera rutan Länka om det infogade grafikobjektet ska ändras så fort någon ändrar originalgrafikfilen.  
Flytta och skala grafikobjektet som du vill.  
Arbeta med en grupp av objekt  
Flera objekt kan markeras tillsammans, grupperas, kombineras, sammansmältas, subtraheras och skäras.  
Gemensam markering har kortast verkan: så fort du klickar på ett annat ställe på sidan upphävs markeringen igen.  
Gruppering och kombination gäller tills du upphäver grupperingen eller kombinationen igen via kommandot på snabbmenyn eller på menyn Ändra.  
Du kan också kombinera de här kommandona, t.ex. sammanfoga flera grupperingar till en enda grupp, lägga till en kombination och sammanfoga resultatet som grupp eller som kombination och så vidare.  
Gruppering av objekt  
Du kan sammanfoga flera objekt till en gruppering.  
Alla ändringar som du sedan gör av grupperingen påverkar alla delobjekt i grupperingen.  
Grupperingar kan också flyttas, roteras m.m. som ett enda objekt.  
Om du till exempel ritar en cykel kan du först konstruera ett hjul som består av däck, fälg, ekrar och nav och sedan gruppera de här objekten.  
Nu är det enkelt att rotera hjulet, kopiera det och flytta kopian.  
Sedan ritar du ramen och resten av cykeln och gör en ny gruppering av detta.  
Då kan du redigera det önskade objektet och sedan lämna grupperingen igen.  
Gå in i grupp  
Du går in i en grupp genom att först markera den (klicka på den eller använd tangentbordet - se vidare längre ner).  
Sedan kan du välja mellan att använda ett (snabb )menykommando eller tangenten F3 eller att dubbelklicka på gruppen för att gå in i den.  
Om du går in i gruppen genom att dubbelklicka är inget objekt i gruppen markerat.  
Lämna grupp  
För att lämna en grupp kan du också välja mellan att använda menykommando eller tangentkombinationen Kommando Ctrl +F3 eller att dubbelklicka utanför alla objekt i gruppen.  
När du lämnar en grupp markeras den, vilket innebär att det är lätt att gå in i gruppen och lämna den igen via tangentbordet.  
Visning av gruppen  
För att gruppen och objekten som den innehåller ska framhävas, visas alla objekt som inte finns i gruppen (alltså även andra grupper) i det nya "spökläget "i bleka färger.  
På så sätt är det lätt att se vilka objekt som är tillgängliga för interaktion och vilka som inte är det, och om du just är i en grupp eller inte.  
Navigering mellan objekt i en grupp (eller på en sida)  
Du kan markera varje objekt i tur och ordning, framåt eller bakåt, i en grupp som du har gått in i med F3 eller på en sida, genom att använda tangenterna Tabb och Skift+Tabb.  
Om du trycker på tangenterna upprepade gånger och kommer till det sista objektet åt ett håll markeras det första objektet igen.  
Sätta samman 3D-objekt  
Du kan koppla samman två 3D-objekt till ett enda objekt, vars konturer är summan av de enskilda objekten.  
Infoga ett 3D-objekt i din presentation eller teckning, t.ex. en kub, med hjälp av utrullningslisten 3D-objekt.  
Infoga ett andra 3D-objekt, t.ex. en kula, som är något större än kuben.  
Klipp ut det andra objektet, d.v.s. kulan, till urklippet med Kommando Ctrl +X.  
Klicka på kuben och tryck på F3.  
Infoga kulan från urklippet med Kommando Ctrl +V.  
Kulen är nu en del av kubens grupp.  
Lämna gruppen, t.ex. med Kommando Ctrl +F3.  
Subtraktioner och snittmängder går inte att göra med 3D-objekt.  
3D-objekt  
Förbinda linjer till ett objekt  
Så skapar du en sluten yta av flera linjer i %PRODUCTNAME Draw eller Impress.  
Via funktionen Förbind är det möjligt att kombinera enskilda linjer till ett ytobjekt.  
Gör som i följande exempel:  
1.  
Linjernas start - och slutpunkter skall ligga nära varandra i de tre hörnorna.  
2.  
Markera alla tre linjerna genom att t.ex. dra upp en rektangel som innesluter alla linjer med urvalsverktyget (pilen längst upp i verktygslisten).  
3.  
Öppna snabbmenyn över de markerade objekten och välj sedan kommandot Förbind.  
4.  
Öppna snabbmenyn igen och välj kommandot Slut objekt.  
5.  
Objektet sluts nu och kan bearbetas som yta.  
Anvisningar för %PRODUCTNAME Draw  
Redigera och gruppera objekt  
Redigera färger och texturer  
Redigera text  
Arbeta med nivåer  
Övrigt  
Rotera objekt  
När du klickar på ett objekt första gången, visas de åtta handtagen som du kan använda om du vill ändra storleken.  
Du kan också ändra objektets placering på sidan genom att dra hela objektet.  
Klicka på ikonen för rotation som du hittar på verktygslisten Effekter i %PRODUCTNAME Draw och direkt på verktygslisten i %PRODUCTNAME Impress.  
Om du rör med musen över handtagen, så kommer muspekaren att visa att du kan rotera objektet genom att dra med musen.  
I mitten av objektet ser du en liten cirkel som visar rotationspunkten.  
Om du drar med musen i handtagen i objektets hörn roteras det runt rotationspunkten.  
Om du däremot drar i handtagen på sidornas mitt så roteras objektet i den tredje dimensionen i förhållande till motstående kant.  
Om du klickar en gång till i objektet ser du de normala åtta handtagen igen.  
Men om du i stället dubbelklickar i objektet förändras de åtta handtagen och du ser en textmarkör i mitten av objektet.  
Du kan nu mata in en text som automatiskt är knuten till objektet.  
Det kan förekomma att enstaka störningar syns på bildskärmen.  
Tryck i så fall på tangentkombinationen Kommando Ctrl +Skift+R för att bygga upp bildskärmen på nytt.  
Omvandla text till 3D  
Om en text är markerad kan du omvandla den till ett tredimensionellt objekt med snabbmenykommandot Omvandla till 3D.  
Det skapade 3D-objektet tar upp utrymmet som du har ritat upp för textramen med musen.  
Den tredimensionella texten kan du rotera fritt.  
Klicka på ikonen Rotera på Effekt-utrullningslisten på verktygslisten.  
Om du klickar innanför begränsningsramen och drar med nertryckt musknapp, roterar objektet runt alla axlar samtidigt.  
Om du klickar på ett av de åtta handtagen och drar med nertryckt musknapp, roterar objektet runt en axel.  
Rotationspunkten, som först visas som en liten cirkel i mitten, kan du flytta med musen.  
Om du sedan roterar objektet, roterar det runt den nya rotationspunkten.  
Öppna fönstret 3D-effekter med ikonen 3D-controller.  
Här tilldelar du 3D-objektet t.ex. en annan belysning.  
Fönstret 3D-effekter beskrivs i %PRODUCTNAME -hjälpen.  
Mata in texter  
Om du vill infoga texter i din teckning, kan du välja mellan att texterna skall visas i "normal" formatering, som t.ex. i ett textdokument, eller om du vill behandla texterna som ett grafikobjekt och t.ex. dra ut, krympa eller rotera dem.  
Dessutom kan du mata in en "normal" text i form av en förklaring, alltså i en ram med en pil.  
Öppna utrullningslisten Text på verktygslisten.  
(Om du har aktiverat stödet för asiatiska språk under Verktyg - Alternativ -Språkinställningar -Språk finns här ikoner som du använder om du vill skriva vertikal text.)  
Normal text  
1.  
En "normal" text infogar du med ikonen Text.  
Klicka på ikonen.  
2.  
Den anger positionen och den maximala bredden på textområdet i dokumentet.  
Den här ramen kan växa nedåt för att all text skall få plats om texten är lång.  
Men ramen kan aldrig bli mindre än själva texten.  
3.  
Mata in texten.  
Du kan markera den med musen, eller genom att hålla ner skifttangenten och använda piltangenterna och sedan ändra t.ex. teckensnitt och teckenstorlek på samma sätt som i textdokument.  
Om du klickar utanför texten i dokumentet lämnar du ordbehandlingsläget.  
Om du därefter klickar en gång i texten markeras den som textobjekt.  
Nu kan du t.ex. flytta och rotera objektet.  
Om du dubbelklickar i texten kan du redigera den igen, t.ex. radera tecken eller sätta teckensnittsattribut.  
Anpassa text till ram  
1.  
Den anger position och storlek för texten som du sedan kan börja mata in direkt.  
2.  
Mata in en text och klicka sedan på ett fritt ställe i dokumentet.  
Den inmatade texten dimensioneras automatiskt till höjd och bredd så att den passar in i ramen.  
Förklaring  
1.  
Med ikonen Förklaring drar du från den punkt på vilken förklaringspilen skall visa till den punkt där förklaringstexten skall stå.  
När du släpper musknappen kan du bearbeta storleken på förklaringsramen.  
2.  
När du vill mata in texten i förklaringen, dubbelklickar du på ramen.  
Den breda gråa kanten på förklaringsramen visar att du nu befinner dig i textbehandlingsläget.  
3.  
Mata in förklaringstexten.  
4.  
Ändra linjens egenskaper genom att klicka på linjen, öppna snabbmenyn och välja Linje.  
Klicka på fliken Linje och välj pilspetsar för linjerna i kombinationsfältet Stil.  
Förse bitmap med text  
Om du t.ex. vill förse en pixelbild i JPEG-format med en text, gör du så här:  
1.  
Öppna ett nytt teckningsdokument.  
2.  
Infoga pixelbilden genom att välja Infoga - Grafik.  
3.  
Upphäv markeringen av den infogade pixelbilden genom att klicka någon annanstans i dokumentet.  
4.  
Öppna utrullningslisten Text på verktygslisten och klicka t.ex. på ikonen Anpassa text till ram.  
5.  
Rita upp en ram på pixelbilden med musen och mata sedan in texten.  
6.  
Du kan markera texten om du vill och ge den en annan teckenfärg.  
Bakgrunden till texten är automatiskt transparent.  
7.  
Markera pixelbilden tillsammans med texten genom att t.ex. rita upp en markeringsram runt båda med musen.  
På statuslisten står då t.ex. "Markerad 2 Ritobjekt".  
8.  
Välj Arkiv - Exportera.  
I dialogrutan Exportera väljer du filtypen "JPEG - Joint Photographic Experts Group" och matar in ett namn.  
Markera rutan Markering så att bara de markerade objekten exporteras.  
9.  
Klicka på Spara.  
I en dialogruta kan du ställa in alternativ för kvaliteten på den skapade JPG-bilden.  
Ju högre kvaliteten är, desto större blir den skapade filen.  
Välkommen till %PRODUCTNAME Draw-hjälpen  
Hjälp till %PRODUCTNAME Draw  
Hjälp till hjälpen  
Menyer  
Här hittar du beskrivningen av alla menyer med undermenyer och dialogerna som kan öppnas.  
Arkiv  
Denna meny innehåller kommandon som du använder när du hanterar dokument i sin helhet.  
Du kan t.ex. skapa ett nytt dokument, öppna, stänga och skriva ut dina dokument, ange dokumentegenskaper med mera.  
När du vill avsluta ditt arbete med %PRODUCTNAME Draw klickar du på menykommandot Avsluta.  
Öppna...  
Spara som...  
Exportera...  
Versioner...  
Egenskaper...  
Skriv ut...  
Skrivarinställning...  
Redigera  
Här hittar du bland annat kommandon för att ångra den senaste åtgärden, kopiera och klistra in via urklippet och för att använda funktionen Sök och ersätt.  
Klistra in innehåll...  
Sök och ersätt...  
Duplicera...  
Tona över...  
Fältkommando...  
Radera sida...  
Radera nivå...  
Länkar...  
Image map  
Hyperlänk  
Visa  
Denna meny kombinerar kommandon som du använder till att styra hur dokumentinnehållet visas på bildskärmen.  
Skala...  
Infoga  
På den här menyn är alla kommandon sammanfattade som används till att infoga nya element i dokumentet, som t.ex. stödlinjer, skannade objekt, grafik, objekt, symboler och andra filer.  
Sida  
Nivå...  
Infoga fångpunkt / -linje...  
Specialtecken...  
Hyperlänk  
Tabell  
Diagram...  
Ram...  
Fil...  
Format  
Här hittar du kommandona för att ställa in objekt - och sidformateringen.  
När du har markerat objekt ändrar sig menyn och visar då särskilda formatkommandon.  
I den här menyn hittar du också funktionerna för hantering av mallar, t.ex. mallkatalogen och Stylist.  
Linje...  
Yta...  
Text...  
Position och storlek...  
Kontrollfält...  
Formulär...  
Dimensionering...  
Förbindelse...  
Tecken...  
Numrering / punktuppställning...  
Stycke...  
Sida...  
Nivå...  
Verktyg  
Menyn Verktyg innehåller kommandon beträffande lingvistik och diverse programalternativ.  
Här startar du rättstavningskontrollen eller synonymordlistan som kan ge dig förslag på alternativa ord.  
Dessutom kan du ställa in utseendet för symbollister och menyer, konfigurera tangentbordet och göra allmänna standardinställningar för programmet.  
Synonymordlista...  
AutoKorrigering...  
Makro...  
Anpassa...  
Symbollister  
Här hittar du en beskrivning av elementen på symbollisterna i ett aktivt teckningsdokument.  
Objektlisten i teckningsvyn  
På den här objektlisten finns det funktioner som du behöver i det aktuella redigeringsläget.  
Linjestil  
Linjebredd  
Linjefärg  
Listrutorna Ytstil / -fyllning  
Verktygslist  
I standardinställningen är verktygslisten placerad till vänster bredvid dokumentet.  
I denna förankringsbara list finns alla de viktigaste redigeringsmöjligheterna.  
Flera av ikonerna är utrullningslister, som i sin tur innehåller fler ikoner.  
Ikonerna med utrullningslister är markerade med små trekanter.  
Alternativlist  
Du kan aktivera alternativlisten under Visa - Symbollister.  
Standardplaceringen är nedanför arbetsytan.  
På den här förankringsbara listen har du tillgång till viktiga alternativ utan att du behöver öppna några dialogrutor.  
Visa raster  
Hjälplinjer vid förflyttning  
Fäst mot raster  
Fäst mot stödlinjer  
Fäst mot sidmarginaler  
Fäst mot objektram  
Fäst mot objektpunkter  
Tillåt snabbredigering  
Bara textområde kan markeras  
Antyd extern grafik  
Konturläge  
Antyd text  
Visa bara fina linjer  
Funktioner i %PRODUCTNAME Draw  
Här hittar du en överblick över några av funktionerna i %PRODUCTNAME Draw, som är modulen för att arbeta med teckningar i %PRODUCTNAME.  
Utforma och publicera vektorgrafik  
%PRODUCTNAME Draw är ett objektorienterat ritprogram för vektorgrafik.  
Objekten kan vara linjer, rektanglar, tredimensionella cylindrar eller andra kroppar och ytor.  
Alla objekt har ett antal egenskaper, som storlek, färg för ytor, färg för inramning, länkade filer, tilldelade funktioner när du klickar på dem med mera.  
Du kan ändra alla egenskaper när som helst.  
Tack vare vektortekniken kan du rotera objekt hur du vill och ändra deras storlek utan att det medför störande trappstegseffekter i kanterna.  
Och eftersom alla objekt hanteras var för sig, kan du flytta och stapla dem på eller under varandra.  
Skapa 3D-objekt  
I %PRODUCTNAME Draw är du inte begränsad till att arbeta med två dimensioner.  
Du kan även skapa kuber, klot, cylindrar och andra 3D-objekt på sidan, rotera dem fritt och till och med belysa varje objekt med en ljuskälla som kan ställas in på många olika sätt.  
I kombination med de fritt definierbara eller fördefinierade färggradienterna kan du i en handvändning utforma iögonfallande sidor för presentationer inom företaget och på Internet.  
Hantera organisationsscheman  
%PRODUCTNAME Draw arbetar objektorienterat.  
Objekt på en sida kan t.ex. vara rektanglar som innehåller text och som är kopplade till varandra.  
Om du flyttar rektanglar på sidan följer förbindelserna med automatiskt.  
Det gör det lätt för dig att rita upp och administrera organisationsscheman för hela företaget eller enskilda avdelningar.  
Detta gör att det är lätt att ta fram tekniska skisser med förklarande text.  
Rita  
Du ritar räta linjer, frihandslinjer, bézierkurvor och alla typer av rätvinkliga och andra figurer på vanligt sätt.  
3D-funktionerna kan användas till att snabbt ta fram 3D-objekt, som t.ex. parallellepipeder, koner, cylindrar, torusar med mera.  
Självklart kan du också rotera dina egna tvådimensionella konturer till den tredje dimensionen.  
Med hjälp av de här effekterna skapar du snygga 3D-objekt för inbjudningskort, broschyrer och visitkort.  
Utnyttja det stora urvalet av clipart som finns i Gallery, oavsett om det rör sig om vektor - eller pixelgrafik, för att lägga till ytterligare element i dina teckningar.  
Exportera  
Med %PRODUCTNAME Draw kan du snabbt och enkelt t.ex. utforma knappar och ikoner för dina webbsidor och exportera dem som GIF, JPG, PNG eller i andra format.  
Konstruera  
Det finns många funktioner som hjälper dig att skapa exakta teckningar.  
Du kan också tillfälligt anpassa nya objekt till de befintliga objektens kanter och punkter.  
Även i teckningen som sådan är det lätt att infoga måttlinjer, som kan ställas in på många olika sätt.  
Integrera  
Naturligtvis kan du också när som helst integrera texter, tabeller, diagram eller formler från de andra programdelarna i %PRODUCTNAME i dina teckningar.  
Så hittar du den här funktionen...  
Rektangel  
Ellips  
Kurva  
Justering  
Placering  
Menyn Arkiv  
Menyn Arkiv - Exportera...  
Menyn Redigera  
Menyn Redigera - Duplicera...  
Skift+F3  
Menyn Redigera - Tona över... (bara i %PRODUCTNAME Draw)  
Menyn Redigera - Radera sida...  
Menyn Redigera - Radera nivÃ¥...  
Menyn Redigera - FÃ¤ltkommando...  
Menyn Visa  
Menyn Visa - Linjaler  
Menyn Visa - Symbollister - Alternativlist  
Menyn Visa - Symbollister - Presentation  
Ikon på objektlisten:  
Presentationslist på / av  
Menyn Visa - Arbetsvy  
Menyn Visa - Visningskvalitet  
Menyn Visa - FÃ¶rhandsvisning visningskvalitet  
Menyn Vy - Arbetsvy - Teckningsvy  
Ikon ovanför den vertikala rullningslisten:  
Teckningsvy  
Menyn Visa - Arbetsvy - Dispositionsvy  
Ikon ovanför den vertikala rullningslisten:  
Dispositionsvy  
Menyn Visa - Arbetsvy - Diabildsvy  
Ikon ovanför den vertikala rullningslisten:  
Diabildsvy  
Menyn Visa - Arbetsvy - Anteckningsvy  
Ikon ovanför den vertikala rullningslisten:  
Anteckningsvy  
Menyn Visa - Arbetsvy - Flygbladsvy  
Ikon ovanför den vertikala rullningslisten:  
Flygbladsvy  
Menyn Bildskärmspresentation - Bildskärmspresentation  
Tangentkombinationen Kommando Ctrl +F2  
Ikon på verktygslisten:  
Bildskärmspresentation  
Ikon ovanför den vertikala rullningslisten:  
Starta bildskärmspresentation  
Menyn Visa - FÃ¶rhandsvisning  
Menyn Visa - Sida  
Ikon på den horisontella rullningslisten:  
Sidvy  
Menyn Visa - Bakgrund  
Ikon på den horisontella rullningslisten:  
Bakgrundsvy  
Menyn Visa - Bakgrund - Teckning  
Menyn Visa - Bakgrund - Titel  
Menyn Visa - Bakgrund - Anteckningar  
Menyn Visa - Bakgrund - Flygblad  
Menyn Visa - Nivå  
Ikon på den horisontella rullningslisten:  
Nivåvy  
Menyn Infoga  
Menyn Infoga - Sida...  
Snabbmeny på flikarna:  
Infoga sida...  
Klicka på det fria området bredvid flikarna  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga sida  
Menyn Infoga - Duplicera sida  
Menyn Infoga - Sidor från disposition  
Menyn Infoga - Översiktssida  
Menyn Infoga - Nivå (bara i %PRODUCTNAME Draw)  
I nivåläge: snabbmenyn på flikarna:  
Infoga nivå...  
Menyn Infoga - Stödpunkt / -linje (bara i %PRODUCTNAME Draw)  
Snabbmeny:  
Infoga stödpunkt / -linje  
Snabbmeny - Redigera stödpunkt / Redigera stödlinje  
Menyn Infoga - Tabell  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga %PRODUCTNAME Calc-tabell  
Menyn Infoga - Fil... (när en fil har valts ut)  
Ikon på utrullningslisten Infoga på verktygslisten  
Fil  
Menyn Infoga - Fältkommando  
Menyn Infoga - Fältkommando - Datum (fast)  
Menyn Infoga - Fältkommando - Datum (variabelt)  
Menyn Infoga - Fältkommando - Klockslag (fast)  
Menyn Infoga - Fältkommando - Klockslag (variabelt)  
Menyn Infoga - Fältkommando - Sidnummer  
Menyn Infoga - Fältkommando - Författare  
Menyn Infoga - Fältkommando - Filnamn  
Menyn Format  
Menyn Format - Dimensionering  
Ikon Måttlinje på utrullningslisten Linjer  
Menyn Format - FÃ¶rbindelse...  
Menyn Format - Sida...  
Menyn Format - Sida... - fliken Sida  
Menyn Format - Sida... - fliken Bakgrund  
Menyn Format - Ã„ndra sidlayout...  
Menyn Visa - Nivå, därefter Ändra nivå... på snabbmenyn  
Menyn Format - Formatmallar - Sidformatmall...  
Menyn Verktyg  
Menyn Verktyg - Avstavning  
Redigera...  
Menyn Bildskärmspresentation  
Menyn BildskÃ¤rmspresentation - DiabildsvÃ¤xling  
Menyn Bildskärmspresentation - Animation  
Menyn Bildskärmspresentation - Effekt  
Ikon på verktygslisten:  
Effekt  
Menyn Bildskärmspresentation - Interaktion...  
Ikon på verktygslisten:  
Interaktion  
Menyn BildskÃ¤rmspresentation - PresentationsinstÃ¤llningar...  
Menyn BildskÃ¤rmspresentation - Individuell bildskÃ¤rmspresentation...  
Menyn Ändra  
Menyn Ändra - Omvandla (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Omvandla - Till kurva (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla - Till kurva (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Omvandla - Till polygon (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla - Till polygon (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Omvandla - Till 3D (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla - Till 3D (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Omvandla - Till 3D-rotationsobjekt (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla - Till 3D rotationsobjekt (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Omvandla - Till bitmap (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla - Till bitmap (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Omvandla - Till Metafil (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla - Till Metafil (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Omvandla - Till kontur (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Omvandla - Till kontur (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Placering - Framför objektet (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Placering - Framför objektet (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Ikon på verktygslisten / placering:  
Framför objektet  
Menyn Ändra - Placering - Bakom objektet (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Placering - Bakom objektet (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Ikon på verktygslisten / placering:  
Bakom objektet  
Menyn Ändra - Placering - Byt (%PRODUCTNAME Draw)  
Snabbmeny vid markerat objekt - Placering - Byt (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Ikon på verktygslisten / placering:  
Byt  
Menyn Ändra - Namnge objekt...  
Snabbmeny till objektet - Namnge objekt...  
Menyn Ändra - Kombinera (%PRODUCTNAME Draw)  
Snabbmeny Kombinera (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Upphäv kombination (%PRODUCTNAME Draw)  
Snabbmeny Upphäv kombination (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Förbind (%PRODUCTNAME Draw)  
Snabbmeny Förbind (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Bryt ner (%PRODUCTNAME Draw)  
Snabbmeny Bryt ner (%PRODUCTNAME Draw och %PRODUCTNAME Impress)  
Menyn Ändra - Former (%PRODUCTNAME Draw)  
Snabbmeny vid markerade objekt Former (%PRODUCTNAME Impress och %PRODUCTNAME Draw)  
Menyn Ändra - Former - Sammansmält (%PRODUCTNAME Draw)  
Snabbmeny vid markerade objekt Former - Sammansmält (%PRODUCTNAME Impress och %PRODUCTNAME Draw)  
Menyn Ändra - Former - Dra ifrån (%PRODUCTNAME Draw)  
Snabbmeny vid markerade objekt Former - Dra ifrån (%PRODUCTNAME Impress und %PRODUCTNAME Draw)  
Menyn Ändra - Former - Skär av (%PRODUCTNAME Draw)  
Snabbmeny vid markerade objekt Former - Skär av (%PRODUCTNAME Impress und %PRODUCTNAME Draw)  
Exportera  
Här exporterar du presentationer och teckningar eller markerade objekt till andra grafikformat.  
Om du väljer "Webbsida" som format skapas filerna med hjälp av en AutoPilot.  
Du kan välja om filerna ska sparas i JPEG - eller GIF-format på en lokal lagringsenhet, på en nätverksenhet eller på en Internet-server (om du har skrivrättigheter där).  
Den här dialogrutan är uppbyggd på samma sätt som dialogrutan Spara som.  
Om du vill exportera en fil i dialogrutan Exportera och klickar på Spara öppnas för många format en filterdialogruta där du kan välja önskade exportalternativ.  
Vilken filterdialogruta som öppnas beror på vilket filformat du valt.  
Följande filterdialogrutor finns:  
HTML-export, JPEG alternativ, SVM / WMF / PICT / MET alternativ, BMP alternativ, GIF alternativ, EPS exportalternativ, PNG alternativ, PBM, PPM, PGM-alternativ..  
Det finns mer information om filter i Information om import - och exportfilter.  
Sida...  
Med det här kommandot öppnar du dialogrutan Ställ in sida, där du bl.a. kan definiera pappersformat och sidbakgrund.  
Där kan du välja om inställningarna som du har gjort ska gälla för alla befintliga och framtida sidor eller bara för den aktuella sidan.  
På så vis kan du t.ex. ge varje sida en annan bakgrund.  
Klicka på önskat alternativ.  
Sida  
Här kan du bestämma sidornas formatering.  
Du kan göra diverse förinställningar, t.ex. vilket pappersformat som används, av numrering och marginalbredd.  
I förinställningarna får nya sidor ett format som passar bildskärmen utan marginaler.  
Pappersformat  
Här väljer Du bland de vanligaste pappersformaten.  
Om Du väljer ett pappersforamt här får Du automatiskt i kombinationsfälten Bredd och Höjd de mått som motsvarar Ditt val.  
Om Du gör egna inmatningar i kombinationsfälten Bredd eller Höjd så ändras formatet i listrutan Pappersformat till Användare.  
Format  
Välj ett fördefinierat pappersformat i listrutan Format, eller ange önskat pappersformat i fälten Bredd och Höjd.  
Bredd  
Här anger Du pappersbredden om Du vill ha en avvikelse från standardformatet.  
Höjd  
Här anger du pappershöjden om du vill ha en höjd som avviker från standardformatet.  
Stående  
Ange i detta alternativfält om dokumentet ska visas eller skrivas ut i stående format (portrait).  
Liggande  
Ange i detta alternativfält om dokumentet ska visas eller skrivas ut i liggande format (landscape).  
Pappersmatning  
Om Din skrivare är utrustad med flera pappersmagasin kan Du här bestämma vilket fack som ska användas.  
Det är nödvändigt att välja pappersmagasin (fack) om Du vill ha ett annat pappersformat från och med den andra sidan.  
Sidmarginaler  
I programmet kan Du ange avståndet mellan skrivtecknen och papperets sidokanter.  
Du kan ändra avståndet i respektive rotationsfält.  
Här kan Du också ange olika måttenheter, som automatiskt räknas om.  
Vänster  
I det här kombinationsfältet kan du definiera storleken på vänstermarginalen.  
Höger  
Här kan du definiera storleken på högermarginalen.  
Uppe  
Här definierar du storleken på den övre marginalen.  
Nere  
Här bestämmer du storleken på den undre marginalen.  
Format  
I den här listrutan definierar du numreringstypen.  
Anpassa objekt till sidformat  
Här kan du definiera om du vill att teckningselementen ska placeras även när pappersformatet byts ut.  
På så sätt bibehålls sidlayouten.  
Vid presentationsobjekt anpassas i sidformatmallen teckensnittets höjd i mallen till layouten.  
På så sätt är det t ex möjligt att avbilda en mall-sidlayout på olika sidformat.  
Bakgrund  
Här väljer du sidornas bakgrunder en och en eller alla samtidigt.  
De tillgängliga kommandona motsvarar de i dialogrutan Yta  
Navigator  
Med det här kommandot sätter du på och stänger av Navigator.  
Med Navigator kan du t.ex. snabbt förflytta dig i ett dokumentet med många diabilder eller snabbt växla mellan laddade dokument.  
Navigator är ett förankringsbart fönster.  
Du öppnar Navigator på bildskärmen när ett dokument är öppet genom att välja Redigera - Navigator, klicka på ikonen på funktionslisten eller trycka på funktionstangenten F5.  
Om Navigator döljer viktig text kan du flytta fönstret genom att placera muspekaren på titellisten och hålla ner musknappen.  
Om du dubbelklickar på titellisten förminskas eller förstoras fönstret.  
Om du vill att Navigator-fönstret ska förankras när du flyttar det så håller du ner Kommando Ctrl -tangenten.  
Liveläge  
Med den här ikonen kan Du aktivera eller inaktivera liveläge under en presentation.  
I liveläge aktiverar Du alla öppnade verktygslister och kan redigera och flytta alla objekt på den aktuella sidan, använda effekter och t o m infoga nya objekt.  
Liveläge  
Penna  
Den här ikonen kan Du endast välja när en presentation körs.  
När Du klickar aktiveras eller inaktiveras en penna på bildskärmen, vilken Du kan göra färgmarkeringar med för att t ex framhäva objekt, stryka under viktiga passager, rita in förbindelser m m.  
Penna  
Första sidan  
Visar första sidan i presentationen som aktuell sida.  
Första sidan  
Förra sidan  
Visar föregående sida i presentationen som aktuell sida.  
Förra sidan  
Nästa sida  
Visar nästa sida i presentationen som aktuell sida.  
Nästa sida  
Sista sidan  
Visar sista sidan i presentationen som aktuell sida.  
Sista sidan  
Draläge  
Sidor och objekt som listas i Navigator kan Du infoga i dokumentet genom att dra med musen.  
Med den här ikonen aktiveras infogningsläget, varvid ikonen visas i en av tre olika vyer.  
Infoga som hyperlänk  
Infoga som länk  
Infoga som kopia  
Infoga som hyperlänk  
Markera det här alternativet på undermenyn om Du vill infoga sidor och objekt, som listas i Navigator, på den aktuella sidan som URL:er.  
Infoga som länk  
Markera det här kommandot på undermenyn om du vill infoga sidor och objekt, som du drar från Navigator till den aktuella sidan, som länkar.  
Detta förutsätter att källsidorna eller -objekten redan har sparats.  
Infoga som kopia  
Om Du markerar det här alternativet infogas sidor och objekt, som Du drar från Navigator, som kopior på den aktuella sidan.  
Befintliga sidor  
I den stora listrutan visas de existerande sidorna.  
Om du dubbelklickar på en sidsymbol visas motsvarande sida.  
Öppnade dokument  
I den här listrutan visas namnen på de dokument som öppnats.  
Om Du vill växla till att visa ett annat öppet dokument i Navigator klickar Du på dokumentnamnet.  
Efter varje dokumentnamn visas inom parentes om dokumentet är aktivt eller inaktivt.  
De aktiva dokumentet väljer Du på menyn Fönster.  
Duplicera  
Med det här kommandot duplicerar du ett markerat objekt.  
Antal kopior  
Här anger du hur många kopior du vill göra av det markerade objektet.  
Uppgifterna som följer gäller alltid den senast infogade kopian.  
Använd värden från markering  
Om du klickar på den här ikonen överförs storleken för det markerade objektet till fälten Förskjutning X-axel och Y-axel.  
På detta sätt uppnår du t.ex. att en kopia av en rektangel som inte har roterats skapas i direkt anslutning till originalet.  
Använd värden från markering  
Placering  
Här väljer du var på sidan som kopian ska infogas.  
X-axel  
I det här rotationsfältet anger du om förflyttningen ska göras till höger eller vänster.  
Med negativa tal placerar du objektet till vänster, med positiva till höger.  
Y-axel  
I det här rotationsfältet anger du om förflyttningen ska göras uppåt eller nedåt.  
Med negativa tal flyttar du objektet uppåt, med positiva nedåt.  
Vinkel  
I detta rotationsfält anger du hur många grader som kopian ska roteras när den infogas.  
Förstoring  
Här kan du välja om kopian ska infogas i originalstorlek eller om den ska förminskas eller förstoras.  
Bredd  
Här anger du den infogade kopians bredd.  
Höjd  
Här anger du den infogade kopians höjd.  
Färger  
När du skapar flera kopior av ett objekt kan du definiera en färggradient från den första till den sista kopian som infogas.  
Start  
Här definierar du vilken färg det först infogade objektet ska ha.  
Slut  
Här definierar du vilken färg det sist infogade objektet ska ha.  
Radera sida  
Med det här kommandot raderar du den aktuella sidan.  
Innan den raderas slutgiltigt måste du bekräfta raderingen.  
Det går bara att välja det här kommandot i teckningsvyn och om presentationen består av flera sidor.  
Radera nivå  
Med det här kommandot raderar du den aktuella nivån.  
Det här kommandot är bara aktivt om du har infogat en nivå.  
Innan nivån raderas slutgiltigt måste du bekräfta raderingen.  
Det går bara att välja den här menypunkten när du har aktiverat nivåvyn.  
Tona över  
Här kan du göra en övergång mellan två markerade, slutna ritobjekt i ett ställbart antal steg.  
%PRODUCTNAME beräknar och ritar mellanstadiernas form och fördelar dem jämnt mellan ursprungsobjekten.  
Den här funktionen är bara tillgänglig när du har markerat två objekt.  
Resultat blir ett nytt gruppobjekt som du kan fortsätta att redigera.  
Inställningar  
Här anger Du inställningar för toningseffekten för två ritobjekt som görs till ett gruppobjekt.  
Steg  
Här kan Du ange det antal steg som ritningsobjekten ska tonas över med.  
Tona över attribut  
Markera det här alternativet om Du vill att objektens attribut (t ex linje - och fyllningsfärg) ska tas med i övertoningen.  
Samma orientering  
Om Du markerar det här alternativet sker övertoningen tvådimensionellt på pappersytan.  
Om alternativet inte är markerat sker en fri rotationen mellan det första och andra objektet.  
Redigera fältkommando  
Här redigerar du formateringen av infogade fältkommandon för datum, klockslag, författare, sidnummer och filnamn.  
Placera textmarkören direkt framför fältkommandot först.  
Fälttyp  
Du kan ändra typ vid behov.  
Fast  
En "fast" fältfunktion fastställer datum eller klockslag när kommandot infogas.  
Variabel  
En "variabel" fältfunktion uppdaterar innehållet varje gång som dokumentvyn uppdateras på bildskärmen.  
Format  
I den här listrutan väljer du formatering för det redigerade fältkommandot.  
Alternativlist  
Med det här kommandot kan du sätta på eller stänga av alternativlisten.  
På alternativlisten har du tillgång till alla alternativ som du ofta behöver när du redigerar %PRODUCTNAME Impress-dokument.  
Linjaler  
Med det här kommandot sätter du på respektive stänger av linjalerna.  
Linjalerna visar positionen för markören och markerade objekt.  
Från linjalerna kan du dra ut stödlinjer på sidan.  
Presentation  
Med det här kommandot öppnar du en liten dialogruta där du kan välja viktiga menykommandon.  
Infoga sida...  
Ändra sidlayout...  
Sidformatmall...  
Teckningsvy  
Med det här kommandot aktiverar du teckningsvyn.  
Dispositionsvy  
Med den här funktionen aktiverar du dispositionsvyn.  
I dispositionsvyn kan du skriva in överskrifterna för de enskilda diabilderna i en presentation.  
Dessutom kan du ordna diabilderna och ändra dispositionsnivån för posterna.  
Det gör du med hjälp av ikonerna Nivå uppåt, Nivå nedåt, Uppåt och Nedåt på textobjektlisten.  
Om du använder tangentbordet kan du ställa markören i början på en rad och trycka på tabbtangenten så flyttas raden en nivå nedåt i hierarkin.  
Om du vill flytta raden en nivå uppåt trycker du dessutom på skifttangenten.  
Om markören inte står i början av en rad, eller om det finns en markering i texten när du trycker på tabbtangenten, infogas bara en tabb på raden utan att dispositionen påverkas.  
Den första dispositionsnivån innehåller de enskilda diabilderna.  
De lägre nivåerna motsvarar överskrifterna till diabilderna.  
Diabildsvy  
Med den här funktionen aktiverar du diabildsvyn.  
I den här vyn kan du visa diabilderna (sidorna) i förminskad storlek, precis som på ett ljusbord.  
Anteckningsvy  
Med den här funktionen aktiverar du anteckningsvyn.  
Texten visas inte vid bildskärmspresentationen.  
Flygbladsvy  
Med den här funktionen aktiverar du flygbladsvyn.  
I flygbladsvyn kan du förminska flera diabilder från en presentation så att de får plats på en sida och sedan skriva ut dem.  
Bildskärmspresentation  
Med det här kommandot startar du en bildskärmspresentation.  
Förinställningarna för en bildskärmspresentation gör du under Bildskärmspresentation - Presentationsinställningar....  
Du kan också starta bildskärmspresentationer genom att klicka med musen på ikonen Starta bildskärmspresentation på symbollisten ovanför den lodräta rullningslisten eller på verktygslisten.  
På snabbmenyn i arbetsområdet hittar du kommandot Bildskärmspresentation, som också utlöser en presentation.  
Du kan även använda kortkommandot Kommando Ctrl +F2.  
Sida  
Med det här kommandot väljer du sidvyn.  
Detta är standardläget när programmet har startats.  
Bakgrund  
Med det här kommandot väljer du bakgrundsvyn.  
I bakgrundsvyn skapar och redigerar du bakgrundselement som inte ska förändras vid presentationen.  
Teckning  
Med det här kommandot kan du välja bakgrundssida till teckningsvyn.  
Rubrik  
Med det här kommandot kan du välja bakgrundssida till rubriksidan.  
Anteckningar  
Med det här kommandot kan du välja bakgrundssida till anteckningsvyn.  
Flygblad  
Med det här kommandot kan du välja bakgrundssida till flygbladsvyn.  
Nivå  
Med det här kommandot väljer du nivåvyn för redigeringen av en sida.  
I nivåvyn kan du flytta och redigera diabildens (sidans) teckningselement på olika nivåer.  
Även om det finns flera nivåer förblir alla teckningselement på de olika nivåerna synliga eftersom varje nivå är transparent.  
Vid behov kan du spärra åtkomsten till en nivå, göra objekten på nivån osynliga och bestämma om en nivå ska kunna skrivas ut.  
Om du vill ändra egenskaperna för en nivå öppnar du dialogrutan Ändra nivå genom att dubbelklicka på fliken till den nivå som du vill ändra.  
Om du bara vill ändra synligheten för alla objekt på en nivå klickar du en gång på fliken för motsvarande nivå samtidigt som du håller ner skifttangenten.  
Nivåns namn visas på ett särskilt sätt (t.ex. i blått eller kursivt) för att antyda att objekten som finns här inte längre är synliga.  
Om du markerar ett objekt ser du i ett fält på statuslisten på vilken nivå det markerade objektet ligger.  
Förhandsvisning  
Med detta kommando kan du se ett förhandsvisningsfönster, som visar hur den aktuella sidan kommer att se ut vid en presentation.  
Vid växling till bakgrundsläget visas förhandsvisningen automatiskt.  
På så sätt kan du kontrollera ändringar snabbare.  
Även om du växlar till dispositionsläget visas förhandsvisningsfönstret.  
Visningskvalitet  
Den här menyn innehåller kommandon som definierar om dokumentet ska visas i färg.  
Den visningskvalitet som du ställer in, sparas automatiskt.  
Färg  
Välj det här alternativet om du har färglagt bakgrunder, text eller andra objekt i en presentation eller en bild och vill att de ska visas i färg.  
Gråskalor  
Välj det här alternativet om du hellre vill se ditt alster i gråskalor.  
Färger visas då som nyanser i grått.  
Intensitet för den gråa färgen varieras beroende på vilken färg som använts.  
Svartvitt  
Om du väljer det här alternativet sker visningen i svartvitt utan färger eller gråskalor.  
En svart skuggning visas t.ex. vit med svart ram.  
Förhandsvisning visningskvalitet  
Med det här kommandot kommer du till en undermeny där du väljer hur många färger som visas i förhandsvisningen.  
Förhandsvisning visningskvalitet är bara tillgänglig om du har aktiverat förhandsvisning.  
Arbetsvy  
Här kan du ställa in önskad arbetsvy.  
I stället för att gå via menyn när du vill växla till respektive läge, kan du klicka på någon av ikonerna som finns uppe i högra kanten av dokumentet.  
Infoga sida  
Med det här kommandot öppnas en dialogruta, där du kan välja vilken mall den nya sidan i dokumentet ska baseras på.  
Namn  
I den här textrutan skriver Du namnet på den nya sidan.  
Välj en AutoLayout  
I den här listrutan kan Du välja önskad layout.  
Nedanför listrutan anges innehållet i den markerade layouten i form av stolpar.  
Visa  
Här kan Du ange om Du vill att en bakgrund med motsvarande objekt ska visas i arbetsområdet.  
Bakgrund  
Markera det här alternativet om den bakgrund som används i layouten ska visas i arbetsområdet.  
Objekt på bakgrunden  
Markera det här alternativet om Du vill att de ritningselement som placerats på bakgrunden ska visas i arbetsområdet.  
Infoga nivå  
Med det här kommandot kan du infoga en teckningsnivå till i det aktuella dokumentet.  
Som standard används bara nivåerna Layout och Controls.  
Vid mer komplicerade teckningar kan du slå samman bestämda teckningselement på en nivå genom att lägga till fler nivåer.  
Det maximala antalet nivåer är begränsat till 65 535.  
Med hjälp av kommandot Visa - Nivå visas de nivåer som finns i dokumentet som flikar, direkt under arbetsområdet.  
Markera en nivå genom att klicka på motsvarande flik.  
Namn  
I detta textfält anger du namnet på den nya nivån.  
Egenskaper  
I det här området väljer du bland alternativen Synlig, Utskrivbar och Spärrad.  
Synlig  
Om den här rutan är markerad visas teckningselementen på den aktuella nivån på bildskärmen.  
Utskrivbar  
Om den här rutan är markerad visas teckningselementen på den aktuella nivån även på utskriften.  
Spärrad  
Om den här rutan är markerad går det inte att markera teckningselementen på den aktuella nivån och det går alltså inte heller att redigera dem.  
Nytt fästobjekt  
Här kan du definiera en stödpunkt eller en vertikal / horisontell stödlinje.  
Stödpunkter eller stödlinjer hjälper dig att justera teckningselement när du ritar.  
De stödpunkter och stödlinjer som infogas kan användas på alla diabilder (sidor) i det aktuella dokumentet, men visas inte vid presentationer eller på utskrifter.  
Du kan även redigera de infogade stödlinjerna och -punkterna (flytta dem med numerisk exakthet eller radera dem).  
Stödpunkter och stödlinjer har "magnetisk" inverkan på objekt som du placerar i närheten av dem med musen.  
Om du placerar ett objekt eller linjalernas nollpunkt i närheten av en stödpunkt eller stödlinje dras objektet / nollpunkten till denna.  
Det gäller även när du skapar ett objekt genom att dra eller klicka med musen.  
Fästområdet ställer du in på menyn Verktyg - Alternativ - Teckning - Raster Verktyg - Alternativ - Presentation - Raster.  
Du kan även dra in stödlinjer från linjalerna till sidan och flytta dem på sidan med musen.  
Du raderar stödlinjer genom att dra tillbaka dem till linjallisten.  
Där kan du redigera eller radera fästobjektet.  
På snabbmenyn kan du välja om stödlinjerna ska synas eller ej genom att markera / avmarkera Stödlinjer synliga.  
På snabbmenyn kan du välja om stödlinjerna ska ligga framför eller bakom andra objekt på sidan med menypunkten Stödlinjer främst.  
Position  
Här kan du ange stödlinjernas eller stödpunkternas placering.  
Du kan när som helst flytta en infogad stödpunkt eller stödlinje med musen.  
X-axel  
Här kan Du ange en horisontell stödlinjes placering eller en stödpunkts X-koordinat.  
Y-axel  
Här anger Du en vertikal stödlinjes placering eller en stödpunkts Y-koordinat.  
Typ  
Här kan Du välja mellan alternativen Punkt, Vertikal och Horisontell.  
Punkt  
Markera det här alternativet om Du vill infoga en stödpunkt.  
Stödpunkten infogas i form av ett streckat kors.  
Vertikal  
Markera det här alternativet om Du vill infoga en vertikal stödlinje.  
Horisontell  
Markera det här alternativet om Du vill infoga en horisontell stödlinje.  
Redigera stödlinje / -punkt  
I fästobjektens snabbmeny kan du flytta eller radera infogade stödlinjer och stödpunkter.  
Dialogrutan är uppbyggd på samma sätt som Nytt fästobjekt.  
Radera  
Med det här kommandot raderar du den aktuella stödpunkten eller stödlinjen.  
Raderingen sker utan någon kontrollfråga.  
Tabell  
Den infogas centrerat.  
Du får tillgång till funktionerna i %PRODUCTNAME Calc för redigering av tabellen.  
Dubbelklicka på tabellen om du vill redigera den igen.  
Klicka en gång på tabellen om du vill flytta den eller ändra storleken.  
Infoga fil  
Med det här kommandot öppnar du en dialogruta, där du kan infoga en presentations-, HTML - eller textfil i dokumentet.  
Du kan lägga in filer från såväl hårddisken som från Internet.  
Om du ska länka in en fil med en URL måste du ange hela URL:en, d.v.s. inklusive file: / / / eller http: / /.  
Den här dialogrutan motsvarar dialogrutan Öppna.  
Välj Filtyp i listrutan och om du vill infoga en text, en webbsida (HTML-dokument) eller ett presentationsdokument.  
Om Du har valt ett presentations - eller HTML-dokument visas dialogrutan Infoga sidor / objekt.  
Här kan Du, i en trädstruktur, välja de sidor eller objekt som Du vill infoga.  
Om Du har valt ett textdokument visas dialogrutan Infoga text.  
Välj textfilen här.  
Efter det att Du har bekräftat Ditt val i dialogrutan enligt ovan, infogas filen eller objektet / objekten i det aktuella dokumentet.  
Infoga sidor / objekt  
I den här dialogrutan infogar du delar av en %PRODUCTNAME Impress - eller HTML-fil i ett presentations - eller teckningsdokument.  
Om du har valt en fil under Infoga - Fil visas den här dialogrutan.  
Om Du inte väljer något av alternativen infogas hela dokumentet.  
Om Du klickar på plustecknet till vänster om filnamnet kan Du välja enskilda sidor eller objekt i %PRODUCTNAME Impress - eller HTML-dokumenten.  
Alla enskilda sidor visas och om det finns inbäddade objekt visas deras namn på en lägre nivå i strukturen.  
Välj de sidor som Du vill infoga.  
Om Du trycker på skifttangenten och Kommando Ctrl kan Du markera flera sidor samtidigt.  
När Du markerat sidorna visas följande fråga i dialogrutan:  
Vill Du anpassa objekten också?  
Klicka på Ja, om Du vill att objekten ska storleksförändras med sidorna.  
Sidor från ett %PRODUCTNAME Impress-dokument läggs till som nya sidor vid den aktuella sidan i dokumentet.  
Visningsområde  
Här väljer Du vad som ska infogas i det aktuella dokumentet.  
Länk  
Markera det här alternativet om Du vill infoga sidorna som länk.  
Då uppdateras det aktuella dokumentet automatiskt när Du öppnar det nästa gång, om ursprungsdokumentet har ändrats.  
Om Du inte markerar det här fältet infogas kopior av sidorna.  
Radera ej använda bakgrundssidor  
Om Du infogar sidor från en presentation eller teckning kan Du här välja om bakgrundssidor i den infogade filen, som inte används, ska tas med i den aktuella filen eller ej.  
Om Du markerar det här alternativet raderas bakgrundssidor, som inte används, från det aktuella dokumentet.  
Infoga text  
Här kan du infoga en textfil (ren ASCII-text, RTF eller HTML) i ett presentationsdokument.  
Du kan även dra upp en textram innan du infogar texten.  
Texten infogas då i den aktuella textramen (den utvidgas nedåt om det behövs - du kan förminska textramen via Format - Position och storlek om den blir för stor.)  
Visningsområde  
Här väljer du vad som ska infogas i det aktuella dokumentet.  
Länk  
Markera den här rutan om du vill infoga sidorna som länk.  
Då uppdateras det aktuella dokumentet automatiskt när du öppnar det nästa gång, om ursprungsdokumentet har ändrats.  
Om du inte markerar den här rutan infogas en kopia av sidorna.  
Duplicera sida  
Med det här kommandot skapar du en kopia av den aktuella sidan.  
Kopian läggs till som ny sida efter den duplicerade sidan.  
Sidor från disposition  
Med det här kommandot skapar du fler sidor från den första dispositionsnivån för den aktuella sidan.  
Den aktuella sidan kan då antingen raderas eller bibehållas.  
Varje dispositionspunkt på första nivån blir en rubrik och dess underordnade punkter blir till disposition för de nya sidorna.  
Den här funktionen är inte tillgänglig i alla lägen.  
Den här funktionen kan endast aktiveras när det finns en disposition på den aktuella sidan.  
De nya sidorna infogas efter den aktuella sidan.  
I en dialogruta får Du frågan "Vill Du radera sidan "sidans namn"?" Om Du bekräftar med Ja att den aktuella sidan ska raderas så bibehålls endast de två nyskapade sidorna.  
Om Du svarar Nej så bibehålls både den aktuella sidan och de båda nya sidorna.  
Översiktssida  
Med det här kommandot skapar du en översiktssida.  
Den innehåller rubrikerna för de enskilda sidorna som disposition på första nivån och utgör därmed ett slags innehållsförteckning.  
Om den första sidan är markerad, sammanfattar kommandot alla sidor.  
Om en annan sida är markerad, sammanfattas alla efterföljande sidor.  
Fältkommando  
Med det här kommandot öppnar du en undermeny där du kan infoga fältkommandon.  
Fältkommandon som används ofta kan du välja direkt på undermenyn.  
Du kan redigera infogade fältkommandon via Redigera - Fältkommando eller via snabbmenyn.  
Datum (fast)  
Det uppdateras inte.  
Du kan ändra formateringen av ett fältkommando genom att placera textmarkören direkt framför fältkommandot och välja kommandot Redigera - Fältkommando.  
Datum (variabelt)  
Med det här kommandot infogar du aktuellt datum som variabel.  
Det uppdateras varje gång som dokumentvyn uppdateras.  
Klockslag (fast)  
Med det här kommandot infogar du aktuellt klockslag som text i dokumentet.  
Det uppdateras inte i fortsättningen.  
Klockslag (variabelt)  
Här kan du infoga aktuellt klockslag som variabel i dokumentet.  
Den uppdateras varje gång dokumentvyn byggs upp igen.  
Sidnummer  
Här infogar du det aktuella sidnumret som fältkommando i dokumentet.  
Formateringen anpassas till den typ som du har ställt in på menyn Format - Sida... i området Numrering.  
Sedan visas aktuellt sidnummer på varje sida.  
Författare  
Här kan du infoga ditt förnamn och efternamn som fältkommando i dokumentet.  
Dessa data hämtas från Verktyg - Alternativ - %PRODUCTNAME - Användardata.  
Filnamn  
Här kan du infoga det aktuella dokumentets filnamn som fältkommando.  
Om du inte har sparat dokumentet ännu är filnamnet tomt.  
Mallkatalog  
Här öppnas en dialogruta, där du kan skapa, ändra och välja mallar.  
Här kan du dessutom administrera de mallar som används i det aktuella dokumentet.  
Alla inställningar i den här dialogrutan hör till de indirekta formateringarna.  
I Stylist har du tillgång till samma funktioner med undantag för administrationen av mallar.  
Malltyp  
%PRODUCTNAME Impress använder som standard malltyperna grafikobjektmallar och presentationsobjektmallar.  
Lista över mallar  
Den mall som används för närvarande är markerad.  
Om du vill välja en annan mall markerar du önskad mall i listrutan.  
På snabbmenyn finns det kommandon, med vilka du kan skapa en ny mall, radera en mall som du har skapat eller ändra den markerade mallen.  
Mallkategori  
För att listan ska bli överskådlig är de färdiga mallarna indelade i flera olika kategorier.  
Välj en annan mallkategori för den aktuella malltypen om den önskade mallen inte visas i listrutan Mallar.  
Alla mallar  
Alla mallar av den aktuella malltypen visas.  
Använda mallar  
Alla mallar av den aktuella malltypen, som används i det aktuella dokumentet, visas.  
Användardefinierade mallar  
Alla mallar av den aktuella malltypen, som definierats av användaren, visas.  
Hierarkiskt  
Mallarna av den aktuella malltypen visas i en hierarkisk struktur.  
Den här vyn liknar katalogstrukuren på en hårddisk.  
Klicka på plustecknet framför mallens namn om Du vill se mallarna på den lägre nivån.  
Nytt...  
Med den här kommandoknappen öppnas dialogrutan Grafikobjektmallar med ett antal flikar.  
Ändra...  
Klicka på den här kommandoknappen om Du vill ändra i den mall som är markerad i listrutan eller kontrollera de aktuella inställningarna för mallen.  
Om Du valt grafikobjektmallar visas dialogrutan Grafikobjektmall som på snabbmenyn Nytt.  
Om Du valt presentationsationsobjektmallar varierar dialogrutans innehåll beroende på den objekttyp som är markerad.  
Beroende på vilken objekttyp Du har valt öppnas dialogrutan för Bakgrund, Bakgrundsobjekt, Rubrik, Underrubrik, Disposition 1 - 9 eller Anteckningar.  
Radera...  
Den markerade mallen raderas efter en säkerhetskontroll.  
Du kan endast radera användardefinierade mallar.  
Förvalta...  
Med den här kommandoknappen öppnar Du dialogrutan Förvalta dokumentmallar.  
Du kan även överföra mallar från andra dokument till det aktuella dokumentet.  
Stylist  
Med Stylist kan du tilldela objekt formatmallar och administrera formatmallar.  
Du kan också skapa nya grafikobjektmallar och ändra deras hierarki.  
Dessutom kan du redigera presentationsobjektmallar här.  
Stylist kommer ihåg vilken typ av mall som du valt i en särskild vy och återställer detta tillstånd så snart du växlar tillbaka till denna vy.  
Det förankringsbara fönstret för Stylist kan du låta vara öppet medan du redigerar dokumentet.  
Ändringar som du gör i formatmallarna påverkar alla sidor som använder dessa mallar.  
Om du vill formatera en presentationssida på ett annat sätt än de andra måste du skapa en ny sidformatmall (masterpage).  
Presentationsobjektmallar  
Presentationsobjektmallar innehåller, beroende av objekttyp, olika typer av information.  
Det kan t.ex. vara använt teckensnitt, teckenstorlek, teckenfärg, uppgifter om styckeindrag och textjustering, information om använda tecken för punktuppställningar, linjetyp, ytfyllning (även för bakgrunden) och skuggor.  
Presentationsobjektmallar  
Grafikobjektmallar  
Grafikobjektmallar innehåller information om mallarnas olika attribut.  
Det kan t.ex. vara använd linjetyp och linjefärg, typ av ytfyllning, skugga, teckensnitt, teckenstorlek och teckenfärg samt uppgifter om styckeindrag och textjustering.  
Grafikobjektmallar  
Tilldelningsläge  
Med hjälp av tilldelningsläget kan du använda den aktuella mallen på ett objekt i arbetsområdet.  
När tilldelningsläget är aktiverat ser muspekaren ut som en färgburk.  
När du vill lämna tilldelningsläget klickar du på ikonen igen.  
Tilldelningsläge  
Så här tilldelar du en ny formatmall i tilldelningsläget:  
Flytta muspekaren till objektet som du vill tilldela den aktuella formatmallen.  
Tryck på vänster musknapp.  
Ny formatmall av markering  
Skapar en ny formatmall med det markerade objektets formatering.  
Du ger den nya formatmallen ett namn i dialogrutan Skapa formatmall som visas automatiskt.  
Ny formatmall av markering  
Uppdatera formatmall  
Formatmallen för det markerade objektet uppdateras med formateringarna för objektet som är markerat i arbetsområdet.  
Uppdateringen påverkar direkt alla teckningselement som använder den här formatmallen.  
Uppdatera formatmall  
Formatmallista / formatmallområde / snabbmenyn Nytt... / Ändra... / Radera...  
Här har du tillgång till samma funktioner som i dialogrutan Format - Formatmallar - Katalog.  
Använda mallar  
I det här fältet ser du vilka mallar som används i dokumentet.  
Använda mallar  
Sidformatmall  
Med hjälp av dialogrutan Sidformatmall kan du välja ut sidformatmallar och tilldela presentationen dem.  
Objekten som ingår i sidformatmallen visas bakom de objekt som redan finns på sidan.  
Sidformatmall  
I listrutan väljer du ut en sidformatmall genom att klicka på den.  
Byt bakgrundssida  
Markera den här rutan om Du vill ersätta bakgrundssidan för alla sidor i dokumentet med den nya sidformatmallen (masterpage).  
Avmarkera rutan om Du bara vill förse den aktuella sidan med en ny sidformatmall.  
Radera ej använda bakgrundssidor  
Markera denna ruta om Du vill ta bort alla bakgrundssidor och presentationslayouter som inte längre används i dokumentet.  
Ladda...  
När Du trycker på knappen visas dialogrutan Ladda sidformatmall.  
Här kan Du välja ut en ny sidformatmall bland de sidformatmallar som finns i systemet.  
Ladda sidformatmall  
Här kan du välja en annan sidformatmall och tilldela presentationen den.  
Kategorier  
Här kan du välja bland mallkategorierna Standard, Sidformat och Presentationsbakgrunder.  
De förinställda alternativen i listrutan Mallar beror på vilken kategori du väljer.  
Mallar  
Här visas en lista över layouterna i den aktuella mallkategorin.  
Tillgängliga alternativ varierar beroende på vad du valt under Kategori.  
Fler>>  
Om du klickar på den här kommandoknappen utökas dialogrutan med följande funktioner.  
Förhandsvisning  
Markera den här rutan om du vill att den presentationslayout du väljer ska visas i förhandsvisningsfältet.  
Förhandsvisningsfält  
Här visas den presentationslayout som du väljer.  
Alla presentationslayouter har inte synligt text - eller bildinnehåll.  
I förhandsvyn visas endast de synliga objekten hos den första diabilden.  
Beskrivning  
Här visas poster med dokumentinformation för de markerade presentationslayouterna.  
Du kan inte ändra förinställningarna här.  
Rubrik  
Här visas mallens rubrik, om sådan finns.  
Tema  
Här visas temat som rubriken hämtats från, om det är tillgängligt.  
Nyckelord  
Eventuella nyckelord som angetts för rubriken visas här.  
Beskrivning  
I tillämpliga fall visas en kort beskrivning av presentationslayouten här.  
Fler<<  
Om du klickar på den här kommandoknappen visas dialogrutan utan tilläggsalternativen.  
Ändra sidlayout  
Här visas en dialogruta där du kan påverka sidans utseende.  
Men textelement kan eventuellt komma att flyttas för att ge plats åt nya grafikobjekt och ramar som tillkommer.  
Namn  
Här anger du önskad beteckning för den nya sidan eller den nya diabilden.  
Standardbeteckningen är Sida X, där X är ett löpnummer.  
AutoLayout  
Klicka på önskad layout i listrutan.  
Nedanför listrutan anges innehållet i den markerade layouten i form av stolpar.  
Visa  
Här kan Du välja vilka element i AutoLayouten som inte ska visas.  
Bakgrund  
Markera det här alternativet om den bakgrund som används i layouten ska visas i arbetsområdet.  
Objekt på bakgrunden  
Aktivera det här fältet om du vill att teckningselementen som placerats på bakgrunden ska visas i arbetsområdet.  
Byta namn på sidan  
Med det här kommandot kan Du byta namn på en befintlig sida eller en bakgrundssida (i presentationslayouten).  
Markera fliken för önskad sida och välj kommandot på snabbmenyn.  
Sedan kan Du skriva in det nya namnet för sidan direkt på sidfliken.  
Presentationsobjektmall för dispositioner  
Här kan du ändra en presentationsobjektmall för en rubrik, underrubrik, disposition eller anteckning.  
Grafikobjektmallar  
Här kan Du skapa en grafikobjektmall.  
Dimensionering  
Förbindelse  
Presentationsobjektmallar  
Här kan Du ändra presentationsobjektmall för en rubrik, underrubrik, disposition eller anteckning.  
Bakgrundsobjekt  
Här kan Du ändra presentationsobjektmallen för ett bakgrundsobjekt.  
Bakgrund  
Här kan Du ändra presentationsobjektmallen för en bakgrund.  
Ändra nivå  
Här kan du ändra några parametrar för sidans aktuella nivå.  
Du kan bestämma om den aktuella nivån ska döljas, spärras och om nivån ska skrivas ut.  
Dialogrutan Ändra nivå öppnar Du med kommandot Ändra nivå... på flikarnas snabbmeny, när Du aktiverat nivåvyn.  
I %PRODUCTNAME Draw (för teckningsdokument) kommer Du även åt menyn via menykommandot Format - Nivå...  
Med Visa - Nivå eller ikonen Nivå vy underst till vänster visar eller döljer Du visningen av flikarna för de olika nivåerna.  
Namn  
Här anger Du en ny beteckning för den aktuella nivån eller accepterar standardnamnet.  
Alternativ  
Med hjälp av kryssrutorna anger Du egenskaperna för den aktuella nivån.  
Synlig  
Markera kryssrutan när ritelementen på den aktuella nivån ska visas på bildskärmen.  
Om innehållet på nivån inte ska synas (t ex egna hjälplinjer för placering i valfria vinklar, kommentarer) så avmarkerar Du rutan.  
Utskrivbar  
Markera denna ruta när ritelementen på den aktuella nivån ska skrivas ut.  
Spärrad  
Markera denna ruta om ritelementen på den aktuella nivån inte längre får markeras, flyttas eller förändras.  
På en spärrad nivå kan Du inte lägga till fler ritelement.  
Byt namn på nivå  
Med detta kommando byter Du namn på en befintlig nivå.  
Markera fliken för motsvarande nivå och välj kommandot på snabbmenyn.  
Därefter skriver Du in det nya nivånamnet direkt på fliken.  
Du kan bara radera och byta namn på nivåer som Du själv har skapat, alltså inte de förinställda nivåerna.  
Dimensionering  
Här definierar du egenskaper för valfria mått, t.ex. mått för objekt.  
Du kan definiera de enskilda attributen och läget för måttet.  
På menyn Format - Linje kan du göra fler inställningar för linjen, linjestilen och linjesluten.  
Dimensioneringen gör du via ikonen Måttlinje på utrullningslisten Linjer på verktygslisten.  
Linje  
I det här området gör du inställningar för dimensioneringen av objekt.  
Du kan ange avståndet mellan dimensioneringslinjerna och objektet, hjälplinjernas längd och önskad visning av dimensioneringen.  
Linjeavstånd  
Här definierar du avståndet mellan dimensioneringslinjen och objektet.  
Hjälplinjeöverhäng  
Här definierar du hur långt hjälplinjerna ska sticka ut utanför dimensioneringslinjen.  
Hjälplinjeavstånd  
Här bestämmer du avståndet mellan hjälplinjerna och objektet.  
Vänster hjälplinje  
Om du vill ändra längden på den vänstra hjälplinjen ställer du in måttet i rotationsfältet.  
Höger hjälplinje  
Om du vill ändra längden på den högra hjälplinjen ställer du in måttet i rotationsfältet.  
Måttlinje nedanför objekt  
Aktivera den här rutan om du vill rotera dimensioneringen 180 grader.  
Etikett  
I det här området definierar du positionen för måttangivelsen i förhållande till dimensioneringslinjen.  
Textposition  
I det här alternativfältet väljer du positionen för måttangivelsen.  
Du har möjlighet att placera visningen av måttet ovanför, genom eller nedanför dimensioneringslinjen.  
Automatiskt vertikal  
Om markerar den här rutan bestäms den optimala vertikala placeringen för måttangivelsen.  
Automatiskt horisontell  
Om du markerar den här rutan så bestäms den optimala horisontala placeringen för måttangivelsen.  
Visa enhet  
Markera det här fältet om du vill att måttenheten för dimensioneringen ska visas.  
Välj en måttenhet i listrutan eller välj "Automatiskt".  
Parallell med hjälplinje  
Med det här alternativet definierar du att dimensioneringen ska placeras parallellt med dimensionseringslinjen.  
Förbindelse  
Här väljer du alla egenskaper för förbindelser.  
Du kan välja linjeförskjutning, linjeavstånd och linjetyp för förbindelser.  
Typ  
Här väljer du typ av förbindelse.  
Du kan välja bland Standardförbindelse, Förbindelselinje, Direktförbindelse och Kurvförbindelse.  
Linjeförskjutning  
Här kan du ange linjeförskjutning i rotationsfälten.  
I förhandsvisningen kan du direkt se effekten av ändringarna.  
Linje 1  
I det här rotationsfältet ställer du in önskad linjeförskjutning för linje 1.  
Linje 2  
I det här rotationsfältet ställer du in önskad linjeförskjutning för linje 2.  
Linje 3  
I det här rotationsfältet ställer du in önskad linjeförskjutning för linje 3.  
Linjeavstånd  
Här kan du ange förbindelsernas linjeavstånd.  
Start horisontellt  
Här anger du hur stort det horisontella linjeavståndet ska vara vid förbindelsens startpunkt.  
Start vertikalt  
Här definierar du hur stort det vertikala linjeavståndet ska vara vid förbindelsens startpunkt.  
Slut horisontellt  
I det här rotationsfältet anger du hur stort det horisontella linjeavståndet ska vara vid förbindelsens slutpunkt.  
Slut vertikalt  
Här definierar du hur stort det vertikala linjeavståndet ska vara vid förbindelsens slutpunkt.  
Du kan förminska och förstora förhandsvisningen genom att klicka med musen.  
Förstora och förminska vyn genom att klicka med den vänstra respektive högra musknappen i förhandsvisningsfönstret.  
Återställ routing  
3 till ursprungsvärdena.  
Placering  
På den här menyn finns kommandona för att lägga grafikobjekt "på varandra".  
Kontroller och andra objekt på kontrollnivån (t ex knappar, kryssrutor osv) i dokumenten ritas alltid upp sist vid bilduppbyggnaden och ligger alltså optiskt sett framför alla andra ritobjekt på sidan.  
Ordningsföljden för markeringar av objekt följer dock fortfarande den interna objektordningen.  
Om Du t ex först ritar en knapp och sedan en rektangel, som delvis täcker knappen, och därefter klickar på det område som de gemensamt upptar på skärmen, så markeras alltid rektangeln.  
Genom att klicka med Alternativ Alt -tangenten nedtryckt markerar Du nästa objekt på samma plats.  
Framför objektet  
Med detta kommando placeras ett objekt framför ett annat objekt.  
Objektet flyttas inte.  
Denna funktion kan du bara använda när minst ett teckningselement är aktiverat.  
Markera det eller de objekt som du vill flytta framåt.  
Välj kommandot.  
Klicka därefter på objektet som ska läggas bakom det markerade objektet eller de markerade objekten.  
Bakom objektet  
Med det här kommandot flyttar du de markerade objekten bakom ett annat objekt.  
Objektet flyttas inte.  
Denna funktion kan du bara använda när minst ett teckningselement är aktiverat.  
Markera det eller de objekt som du vill flytta bakåt.  
Välj kommandot.  
Klicka därefter på objektet som ska läggas ovanpå det markerade objektet eller de markerade objekten.  
Eftersom hänsyn tas till den aktuella ordningsföljden för alla objekt kan detta även leda till en synlig ändring om ett objekt placeras framför eller bakom ett annat objekt även om de båda objekten inte helt eller delvis sammanfaller.  
Objektet, vars position har ändrats i stapeln av objekt, kan placeras ovanpå eller under ett tredje objekt.  
Byt  
Med det här kommandot byter du ordning på objekt.  
Markerade objekt staplas i omvänd ordning.  
Den här funktionen är bara tillgänglig om du har markerat minst två teckningselement samtidigt.  
Mallar  
Här finns kommandon för hantering av mallar.  
Katalog...  
Sidformatmall...  
Avstavning  
Här kan du aktivera eller stänga av avstavningen för textobjekt.  
Avstavningen kan aktiveras eller stängas av styckevis.  
Diabildsväxling  
Här väljer du toningseffekter och hur snabbt diabilderna ska växla för den aktuella sidan eller för de markerade sidorna.  
Effekter  
Med den här kommandoknappen väljer du bland de tillgängliga effekterna för diabildsväxling.  
Effekter  
Effekter  
Här väljer du en effekt för toning mellan sidor (diabilder).  
Hastighet  
I listrutan anger du hastigheten med vilken diabilderna ska växla.  
Du kan välja mellan långsamt, medel eller snabbt.  
Extra  
Med denna kommandoknapp väljer Du bland tillgängliga verktyg för diabildsväxling.  
Välj mellan automatisk och manuell diabildsväxling och om diabildsväxlingen ska ackompanjeras av ljud.  
Verktyg  
Växling  
Här väljer du mellan automatisk, halvautomatisk och manuell diaväxling.  
I dialogrutan Diabildsväxling kan du också välja en ljudfil.  
Diaväxling automatiskt  
Om Du vill ha en automatisk växling mellan de enskilda sidorna (diabilderna), aktiverar Du denna kommandoknapp.  
Diabilden växlas efter att den tid som angetts i rotationsfältet Diavisningstid har förflutit.  
Diaväxling automatiskt  
Halvautomatisk diaväxling  
Välj denna ikon om objekteffekterna ska utföras automatiskt, men sidbytet manuellt.  
Halvautomatisk diaväxling  
Diaväxling manuellt  
Om Du väljer kommandoknappen Diaväxling manuellt sker en växling mellan de enskilda diabilderna först efter det att Du bekräftar detta.  
Diaväxling manuellt  
Visningstid dia  
Här anger Du den tidsrymd efter vilken sidvyn (diabilderna) ska växla.  
Detta fält är bara aktivt om Du valt automatisk växling.  
Ljud  
Aktivera ikonkommandoknappen om en viss ljudfil ska spelas upp vid diabildsväxling.  
Om du klickat på Sök visas standarddialogrutan för val av fil, där du kan välja en ljudfil.  
Ljud  
Sök...  
Med denna kommandoknapp öppnar du dialogrutan Öppna, med vilken du kan ladda en ljudfil.  
Dialogrutan är uppbyggd på samma sätt som Öppna.  
Dessutom finns kommandoknappen Spela upp här.  
Sök...  
Ljudnamn  
I den här listrutan skriver du in namnet på en ljudfil eller väljer en ljudfil i listrutan.  
Uppdatera  
När du har aktiverat den här ikonen visar dialogrutan Diabildsväxling de aktuella inställningarna för en diabild när du har klickat på diabilden.  
Uppdatera  
Tilldela  
Om du vill tilldela en diabildsväxling de valda inställningarna, klickar du här.  
Tilldela  
Förhandsvisning  
Klicka på den här kommandoknappen om du vill se en förhandsvisning av den toningseffekt som du har valt.  
Förhandsvisning  
Animation  
Här styr du sammanställningen och bildföljden för animationssekvensen.  
För att kunna bygga upp en animation behöver du alla objekt som var och är en enskild bild i animationen.  
Du kan växla fram och tillbaka mellan teckningen och dialogrutan, utan att behöva lämna dialogrutan.  
Du kan även infoga animationen i textdokument via urklippet.  
Animation  
När du övertar ett objekt från din teckning, visas det övertagna objektet här.  
När du klickar på kommandoknappen Spela upp ser du animationens förlopp här.  
Med den här ikonen kommer du till den första bilden i din animation.  
Första bilden  
Med den här ikonen kommer du till föregående bild.  
Bakåt  
Med den här ikonen stoppar du animationen.  
Stopp  
Här startas animationen.  
Spela upp  
Med den här ikonen kommer du till den sista bilden i animationen.  
Sista bilden  
Bildnummer  
Här visas den aktuella bildens nummer.  
Om en annan bild ska visas i förhandsvisningsområdet matar du in bildnumret direkt eller ställer in det med pilknapparna bredvid textfältet.  
Visningstid  
I det här rotationsfältet kan du ange den aktuella bildens visningstid.  
Det här fältet är bara aktivt när du har valt alternativet Bitmapobjekt i området Animationsgrupp.  
Mata in tiden direkt, eller ställ in den med pilknapparna bredvid textfältet.  
Visningsförloppet anges i Animator på objektlisten.  
Antal omgångar  
Här kan du ange antal omgångar för animerade bitmapobjekt.  
Posten Max. står för obegränsat antal omgångar.  
Bild  
I det här området hittar du de funktioner som är nödvändiga när du skapar en animation.  
Överta objekt  
Om du vill överta alla markerade objekt i animationen klickar du här.  
De enskilda objekten sammanfogas till en bild.  
Överta objekt  
Överta objekt ett och ett  
Om du vill överta objekten som du har valt till animationen ett och ett, klickar du på den här ikonen.  
Du får en samling bilder som motsvarar antalet objekt som du har markerat.  
Summan för bilderna visas i textfältet Antal.  
Om ett gruppobjekt är markerat övertas även dess enskilda objekt ett och ett.  
Använd den här ikonen om du vill överföra ett markerat animationsobjekt eller en animerad GIF-bild, som infogats på en presentationssida, för att redigera den.  
Vid animerade GIF-bilder kan du redigera de enskilda bildernas visningstid direkt i fönstret Animation.  
Överta objekt ett och ett  
Radera aktuell bild  
Klicka här om du vill radera den aktuella bilden som visas i förhandsvisningsområdet.  
Radera aktuell bild  
Radera alla bilder  
Klicka här om du vill att alla överförda objekt (bilder) ska raderas i animationen.  
Radera alla bilder  
Antal  
Här visas antalet bilder i animationen.  
Animationsgrupp  
I det här området gör du diverse inställningar för animeringsgruppen.  
Du bestämmer hur objekten ska sammanfogas och deras transparensfärg och justering.  
Gruppobjekt  
Markera det här alternativfältet om du vill sammanfoga de enskilda objekten i animationen till ett gruppobjekt.  
Bitmapobjekt  
Om du vill sammanfoga de enskilda objekten i animationen till ett bitmapobjekt, aktiverar du det här alternativfältet.  
Transparensfärg  
I den här listrutan kan du välja en transparensfärg för animationen från den aktuella färgtabellen.  
Men detta är bara möjligt om objekten har sammanfogats till ett bitmapobjekt.  
Anpassning  
Här definierar du de enskilda bildernas justering i förhållande till varandra.  
Alla objekt placeras centrerat som standard.  
Välj justering i listan.  
Skapa  
Välj den här kommandoknappen för att foga in den aktuella versionen av animationen i presentationens diabild.  
Effekt  
Här definierar du en effekt för visningen ett rörligt objekt  
Effekter  
Med den här kommandoknappen väljer du en effekt för det markerade objektet.  
Effekter  
Effekter  
Här väljer du en effekt.  
Om du vill använda effekten Övriga / Flytta längs kurva kan du rita en kurva på diabilden, sedan markera objektet och kurvan samtidigt (håll ner skifttangenten när du markerar) och sedan välja den här effekten.  
Objektets mittpunkt följer kurvan från början till slut.  
Effekterna i området Favoriter har även en ljudeffekt.  
Om du inte vill använda det här ljudet finns samma effekter i de andra områdena där du har möjlighet att avstå från ljud eller tilldela ett valfritt ljud.  
Hastighet  
I den här listrutan definierar du hastigheten för effekten.  
Texteffekter  
Med den här kommandoknappen väljer du texteffekter.  
Texteffekter  
Texteffekter  
Välj en texteffekt.  
Extra  
Med den här kommandoknappen väljer du extraalternativ.  
Extra  
Extra  
Gör objekt osynligt  
Klicka här om du vill att objektet ska bli osynligt efter effekten.  
Gör objekt osynligt  
Tona bort objekt med färg  
Klicka här om du vill tona bort ett objekt med färg.  
Tona bort objekt med färg  
Toningsfärg  
I den här listrutan väljer du en toningsfärg.  
Ljud  
Klicka på ikonen om du vill att en ljudfil ska spelas upp vid diabildsväxlingen.  
Med Sök öppnar du en dialogruta där du kan välja en ljudfil.  
De format som stöds är: .au / .snd (SUN / NeXT Audio), .wav (MS Windows Audio), .voc (Creative Labs (=Soundblaster) Audio), .aiff (SGI / Apple Audio), .iff (Amiga Audio).  
I Windows stöds filformatet WAV.  
Ljud  
Spela upp ljud fullständigt  
Klicka här om Du vill att hela ljudfilen ska spelas upp.  
I Unix spelas alltid hela ljudfilen upp.  
Spela upp ljud fullständigt  
Sök...  
Med den här kommandoknappen öppnar Du dialogrutan Öppna, där Du kan ladda en ljudfil.  
Dialogrutan liknar Öppna.  
Dessutom har Du tillgång till kommandoknappen Spela upp.  
Sök...  
Ljudnamn  
I det här kombinationsfältet väljer du namnet på en ljudfil.  
Ordning  
Klicka på den här kommandoknappen så öppnas en dialogruta, där Du kan definiera i vilken ordningsföljd objekten ska visas.  
Ordning  
Ordningsföljd  
Här definierar du ordningsföljden för presentationen med dra-och-släpp.  
Uppdatera  
Klicka här om Du vill att alla aktuella alternativ som har valts för det markerade objektet ska visas i dialogrutan.  
Uppdatera  
Tilldela  
Om Du vill tilldela det markerade objektet de aktuella inställningarna i dialogrutan, klickar Du här.  
Tilldela  
Förhandsgranskning  
Klicka på den här kommandoknappen så öppnas ytterligare ett fönster med förhandsvisning av den effekt som Du har valt.  
Förhandsgranskning  
Dialogrutans innehåll ändras beroende på vilket alternativ du väljer.  
Åtgärd vid musklick  
Du kan även tilldela åtgärder till grupperade objekt och objekt i 3D-scener.  
Ingen åtgärd  
Välj det här alternativet om Du inte vill utföra någon åtgärd genom att klicka med musen.  
Hoppa till föregående sida  
Om Du väljer det här alternativet sker ett hopp till föregående sida.  
Hoppa till nästa sida  
Om Du väljer det här alternativet sker ett hopp till nästa sida.  
Hoppa till första sidan  
Om Du väljer det här alternativet sker ett hopp till första sidan.  
Hoppa till sista sidan  
Om Du väljer det här alternativet sker ett hopp till sista sidan.  
Hoppa till sida eller objekt  
Om Du klickar med musen på det markerade objektet sker ett hopp till en definierad sida i dokumentet, eller också utförs en åtgärd som är knuten till ett objekt.  
Sida / objekt  
Här visas en lista över alternativen Flygblad, Standard (Flygblad), Standard, Standard (Anteckningar), befintliga Sidor och Sidor (Anteckningar).  
Sida / objekt  
I den här textrutan visas som standard det alternativ Du valt i listrutan Sida / objekt.  
Sök  
Med den här kommandoknappen startar Du en sökning.  
Hoppa till dokument  
När Du valt det här alternativet visas området Dokument.  
Dokument  
Om Du klickar på det markerade objektet laddas ett definierat dokument och den presentationen som ingår i det startas.  
Dokument  
Här kan Du ange namnet för det dokument som ska laddas och vars presentation ska startas.  
Genomsök...  
Dialogrutan Öppna är uppbyggd på samma sätt som Arkiv - Öppna.  
Gör objekt osynligt  
Om Du väljer det här alternativet görs objektet osynligt när Du klickar.  
Spela upp ljud  
Om Du väljer alternativet Spela upp ljud visas rutan Ljud.  
Ljud  
Om Du klickar på det markerade objektet spelas den ljudfil som Du har valt upp.  
Ljud  
Här kan Du ange namnet för den ljudfil som ska laddas och spelas upp.  
Genomsök...  
I den här dialogrutan kan du även välja att det valda ljudet ska spelas upp innan du väljer det som interaktion.  
Om inga ljudfiler installerades när Du installerade %PRODUCTNAME kan Du när som helst installera ljudfilerna i efterhand genom att köra installationsprogrammet och välja alternativet Ändra installation.  
Spela upp  
Klicka på Spela upp om Du vill spela upp ljudfilen.  
Dölj objekt  
Om Du klickar på det markerade objektet döljs det.  
Effekt  
I kombinationsrutan väljer du effekter som ska uppnås när objektet döljs.  
Långsamt  
Klicka här om du vill att objektet ska döljas långsamt.  
Medel  
Aktivera det här alternativfältet om objektet ska döljas i normal hastighet.  
Snabbt  
Klicka här om du vill att objektet ska döljas snabbt.  
Ljud  
I det här omådet väljer du om en ljudfil ska spelas upp.  
Tona ut med ljud  
Klicka här om du vill att en ljudfil ska spelas upp när objektet tonas ut.  
Ljud  
I det här fältet kan du ange namn och sökväg för en ljudfil eller klicka på Genomsök och välj en ljudfil i dialogrutan.  
Spela upp fullständigt  
I Unix spelas alltid hela ljudfilen upp.  
Genomsök...  
I den här dialogrutan kan du även spela upp den valda ljudfilen innan du väljer den som interaktion.  
Vid en standardinstallation av %PRODUCTNAME installeras inga ljudfiler.  
På installation-CD:n finns en katalog med ljudfiler som Du kan installera i efterhand om Du så önskar.  
Spela upp  
Klicka här om Du vill att den valda ljudfilen ska spelas upp.  
Utför program  
I textrutan Program kan Du ange programmets namn.  
Program  
Program  
Här kan du ange namnet på det program som ska laddas och startas.  
Genomsök...  
Dialogrutan är uppbyggd på samma sätt som Arkiv - Öppna.  
Utför makro  
Här kan Du ange ett makro, som ska köras när Du klickar på objektet.  
I textrutan Makro kan Du ange ett makronamn eller också kan Du välja ett makro med kommandoknappen Genomsök....  
Makro  
I det här området finns textfältet Makro och kommandoknappen Genomsök.  
Makro  
Här kan du ange namnet på det makro som ska laddas och startas.  
Genomsök...  
Med den här kommandoknappen öppnar Du dialogrutan Makro, där Du kan välja ett makro.  
Avsluta presentation  
Om du väljer det här alternativet avslutas presentationen när du klickar med musen.  
Presentationsinställningar  
Med det här kommandot öppnar du dialogrutan Bildskärmspresentation.  
Här bestämmer du vilken diabild som ska inleda presentationen och andra alternativ för presentationen.  
Omfång  
Här kan du ange vad presentationen ska omfatta.  
Alla diabilder  
Om du aktiverar det här alternativfältet visas alla diabilder i det aktuella dokumentet i presentationen.  
Från diabild  
Om du inte vill att presentationen ska inledas med första diabilden i det aktuella dokumentet klickar du här.  
I listrutan väljer du den diabild som ska inleda presentationen.  
Individuell presentation  
Om du tidigare har definierat en särskild ordningsföljd för diabilderna i en presentation under Individuell bildskärmspresentation kan du välja den här och köra den som aktuell presentation.  
Typ  
Här anger du i vilket läge (t.ex. helskärm) som presentationen ska köras.  
Standard  
Standardläget är helskärm, där du styr presentationen till sista sidan.  
Den svarta slutsidan innehåller bara en uppmaning att avsluta presentationen genom att klicka med musen.  
Du kan även trycka på valfri tangent.  
Fönster  
Om du väljer det här alternativfältet körs presentationen i dokumentfönstret och inte i helskärm.  
Om du har infogat presentationen som ram, t.ex. i ett textdokument, körs den också i ramen där.  
Om dokumentet ändras i en annan vy medan en presentation körs i ett fönster kan det leda till inkonsekvenser mellan de båda vyerna.  
Om Du t ex raderar ett objekt i dokumentet så kan det hända att objektet ändå visas i presentationen eftersom bitmapmönstret för presentationen redan beräknats i förväg.  
Auto  
I autoläge sker en helskärmsvisning, som upprepas ända tills Du avslutar den.  
Du kan avsluta den automatiska presentationen genom att trycka på Esc-tangenten.  
I det tillhörande rotationsfältet kan Du ange, i sekunder, under hur lång tid en paussida ska visas mellan presentationspassen.  
Efter den angivna paustiden startar presentationen om från början igen.  
Paustid  
Här ställer Du in paustiden mellan upprepningarna av presentationen i autoläge.  
Om värdet är noll visas inte någon paussida.  
Visa logotyp  
Om Du markerar det här alternativet visas %PRODUCTNAME -logotypen på paussidan i autoläge.  
Alternativ  
Medan en presentation pågår visas diabilderna normalt i helskärm.  
Med följande alternativ kan du bestämma hur presentationen ska genomföras.  
När presentationen har startats växlar %PRODUCTNAME Impress automatiskt mellan diabilderna och återgår till normalvy efter den sista diabilden.  
Om du vill avbryta en presentation trycker du på Esc - tangenten.  
Manuell diabildsväxling  
Du växlar till nästa diabild genom att trycka på returtangenten eller högerpilstangenten.  
Du går vidare till nästa animationseffekt på en bild med vänstra musknappen.  
Om Du vill visa föregående diabild trycker Du på vänsterpilstangenten.  
Visa muspekare  
Om Du vill att muspekaren ska synas under presentationen klickar Du här.  
Det här alternativet kan vara lämpligt om Du vill kunna ändra presentationsförloppet genom att välja vissa ritningselement.  
Du kan dessutom använda musknappen för att växla till nästa diabild.  
Muspekare som penna  
Du kan använda muspekaren som penna under presentationen för att markera intressanta områden på bildskärmen.  
Du markerar ett område genom att placera muspekaren på önskat ställe och rita en linje med musknappen nedtryckt.  
Markeringar som Du gör under presentationen sparas inte på diabilderna.  
Det går inte att ändra pennans färg.  
Navigator synlig  
Markera det här alternativet om Du vill att Navigator ska synas under presentationen.  
Tillåt animationer  
Om du markerar det här alternativet kan animerade GIF-objekt och texter visas som animationer.  
I annat fall visas bara första rutan av en animerad GIF-bild eller början på den animerade texten utan animation.  
Diabildsväxling vid musklick på bakgrunden  
Markera det här alternativet om Du vill kunna växla till nästa diabild genom att klicka på bakgrunden.  
Presentation alltid i förgrunden  
Markera det här alternativet om presentationen alltid ska ligga kvar i förgrunden.  
Du behöver då inte bekymra Dig för att andra applikationer (t ex systemmeddelanden eller påminnelser) ska lägga sig framför diabilderna inför all publik.  
Om Du valt fönstervisning för presentationen är det här alternativet inte tillgängligt.  
Individuell bildskärmspresentation  
Med det här kommandot definierar och startar du en presentation, som du har sammanställt av diabilderna i den aktuella presentationen.  
Du kan definiera ett valfritt antal individuella presentationer och ge dem namn.  
De sparas automatiskt i det aktuella dokumentet.  
Presentationens( ernas) namn  
I listrutan visas namnen på de individuella presentationerna.  
Klicka på Ny... om du vill skapa en ny individuell presentation.  
Om du har skapat minst en ny individuell presentation kan du klicka på presentationen i listrutan och sedan köra den.  
Om du vill köra en individuell presentation markerar du den i den stora listrutan.  
Markera dessutom alternativet Använd individuell bildskärmspresentation och klicka på Starta.  
Använd individuell bildskärmspresentation  
Markera den här rutan om den individuella presentation ska visas när du klickat på Starta.  
I annat fall visas hela presentationen i oförändrat skick.  
Ny...  
Redigera...  
Klicka här för att öppna dialogrutan Definiera individuell bildskärmspresentation där du kan redigera den markerade individuella presentationen.  
Kopiera  
Här kan du kopiera den markerade individuella presentationen inom den stora listrutan.  
Den får automatiskt ett namn som du kan ändra - liksom hela den nya presentation - om du klickar på Redigera....  
Starta  
Klicka här för att starta presentationen.  
I annat fall körs hela presentationen.  
Definiera individuell bildskärmspresentation  
Här anger du hur diabilderna ska sättas samman för den individuella presentationen.  
Använd kommandoknapparna >> och << för att sätta samman den individuella presentationen.  
För att ta med en bild klickar Du på >>.  
Klicka sedan på <<.  
Namn  
I detta textfält kan Du ändra namnet på den individuella presentationen.  
Presentationens sidor  
I den vänstra listrutan ser Du den aktuella presentationens diabilder i den ursprungliga ordningsföljden.  
Individuell presentation  
I den högra listrutan ser Du diabildernas ordningsföljd i den individuella presentationen.  
Omvandla  
Här öppnar du en undermeny där du kan omvandla det markerade objektet.  
Till kurva  
De markerade objekten omvandlas till Bézierkurvor.  
Till polygon  
Här omvandlar du objektet till en polygon.  
Genom omvandlingen ändras inte linjernas aktuella utseende.  
De mycket omfattande ändringarna av linjernas uppbyggnad syns först vid redigeringen av punkterna.  
Hela kurvan består efter omvandlingen av ett stort antal raka linjedelar.  
Följande dialogruta visas bara när Du omvandlar en bitmap (pixelgrafik) till en polygon (vektorgrafik).  
Omvandla till polygon  
Förutom att Du kan göra olika inställningar i den här dialogrutan kan Du också förhandsgranska resultatet.  
Inställningar  
I detta område finns inställningsalternativ för omvandlingen.  
Antal färger:  
%PRODUCTNAME Draw skapar en metafil av en bild som består av polygoner.  
Här kan Du ställa in det maximala antalet färgnivåer.  
Punktreduktion:  
Vid inställningen "0 Pixel" skapas alla polygoner.  
Om Du anger ett tal kommer polygoner, som omges av en rektangel med lägre antal pixlar, inte att skapas.  
Fyll hål  
Det händer att färgnivåer inte ligger tillräckligt nära varandra.  
Då kan Du med det här alternativet aktivera en bakgrundsfyllning.  
Fyllningen består av rektanglar vars storlek Du ställer in under Kakelstorlek.  
Kakelstorlek:  
Här ställer Du in storleken för rektanglarna som används för bakgrundsfyllning för alternativet Fyll hål.  
Originalbild:  
Originalbilden (bitmap) som Du har markerat visas i fönstret.  
Vektoriserad bild:  
Med hjälp av knappen Förhandsvisning kan Du se resultatet av Dina inställningar i det här fönstret.  
Framsteg  
Här visas hur konverteringen fortskrider.  
Förhandsvisning  
Här klickar du om du vill se en förhandsvisning.  
Till 3D  
Här omvandlar du objektet till en tredimensionell visning.  
Markeringen omvandlas till en kontur.  
Hänsyn tas då även till linjegeometrierna.  
Exempelvis omvandlas en inramning också till ett 3D-objekt.  
Om du har markerat flera 2D-objekt samtidigt och omvandlar dem till 3D så blir resultatet ett enda 3D-objekt, "scenen".  
Du kan redigera scenen via menyn Ändra - Gå in i gruppering Format - Grupp - Gå in i eller med F3.  
Du kan t.ex. också tilldela dessa objekt en annan färg.  
Enklast lämnar du scenen genom att klicka på ikonen Lämna alla grupperingar på alternativlisten.  
Förutom grupperingar kan Du också omvandla bitmapsbilder och metafilsbilder direkt till 3D-objekt.  
Bitmapsbilder läggs då som textur på ett rektangulärt objekt av motsvarande storlek och omvandlas därefter.  
Detta skiljer sig från en metafil som först upplöses i en grupp av polygoner och för att sedan omvandlas.  
Vid en samtidig omvandling av flera objekt kommer den djupsortering som råder vid 2D-presentationen att användas som information för att skapa 3D-objekt på olika nivåer.  
Då behålls den synlighet som gäller 2D-presentationen.  
Även komplexa Clipart-objekt omvandlas i en förhållandevis snabb process.  
Om ritobjekten innehåller text omvandlas de så att texten fortfarande syns.  
Möjligheterna att utforma objekt är nästan obegränsade.  
Experimentera med verktygen, använd ljuseffekterna, förvrängningseffekterna, texturerna, alternativen som finns i 3D-effekt -fönstret och så vidare.  
Till 3D-rotationsobjekt  
Här omvandlar du objektet till ett tredimensionellt rotationsobjekt.  
Till bitmap  
Här omvandlar du objektet till ett bitmapobjekt (pixelgrafik, rastergrafik).  
I ordlistan hittar du information om bitmap-formatet.  
Denna funktion är detsamma som om Du skulle klippa ut objektet till Urklipp och sedan infoga det igen som en bitmap (med menykommandot Redigera - Infoga innehåll...)  
Till metafil  
Med det här kommandot omvandlar du objektet till ett metafilobjekt (vektorgrafik).  
En kort beskrivning av metafilformatet hittar du i ordlistan.  
Denna funktion är detsamma som om du skulle klippa ut objektet till urklippet och sedan infoga det igen som en metafil (med menykommandot Redigera - Infoga innehåll...)  
Till kontur  
Med det här kommandot omvandlar du det markerade objektet till en grupp av polygoner, som innehåller den kompletta visningsgeometrin för objektet.  
Vid omvandling till kontur tas hänsyn till objektet som sådant, eventuellt teckensnitt i objektet och linjernas geometri med linjestil och pilspetsar.  
På så sätt kan en godtycklig pil skapas, som sedan kan omvandlas till kontur och vidarebearbetas.  
Namn  
Här visas dialogrutan Namn där du kan namnge objektet.  
Namnet som du valt för objektet visas i Navigator och på statuslisten när objektet markerats.  
Det är bara OLE-objekt, grupperade och importerade objekt som kan tilldelas ett namn.  
Vid andra objekt är det här kommandot inte aktivt.  
Namn  
I detta textfält ger Du objektet ett namn.  
Kombinera  
Med det här kommandot skapar du ett nytt teckningselement av de markerade teckningselementen.  
Beroende på de markerade teckningselementens placering i förhållande till varandra skapas nya objektkonturer och eventuellt luckor i objektytan.  
Vidare omvandlas alla teckningselement till Bézierkurvor genom denna kombination.  
Upphäv kombination  
Med det här kommandot kan du dela upp ett teckningselement, som du har skapat med kombinationsfunktionen, i sina enskilda beståndsdelar.  
Teckningselement som du skapar på det här sättet föreligger som Bézierkurvor och får det kombinerade objektets attribut.  
Förbind  
Med det här kommandot skapar du ett nytt linjeobjekt eller en ny Bézierkurva av markerade linjer, delar av linjer eller Bézierkurvor.  
Om inte objekten som ska förbindas har kontakt med varandra skapas en extra förbindelselinje mellan de enskilda linjesegmenten.  
Bryt ner  
Med det här kommandot bryter du ner konturlinjer som är förbundna med varandra.  
Slutna konturlinjer (polygonkurvor, Bézierkurvor) av fyllda teckningselement bryts ner i flera enkellinjer och / eller Bézierkurvdelar.  
Eftersom kurvan inte är sluten efter nedbrytningen kan du inte längre använda ytfyllning.  
Här har du möjlighet att avbryta processen.  
Former  
Här öppnar du en undermeny där du kan använda en mängdoperation på de markerade polygonerna.  
Markera polygonerna gemensamt och välj detta kommando, som Du hittar i markeringens snabbmeny och i %PRODUCTNAME Draw i menyn Ändra.  
Polygonerna sammanfogas till en ny polygon.  
Denna nya polygon får samma attribut som markeringens första (bakersta) polygon.  
Sammansmält  
De markerade polygonerna smälts samman (logiskt ELLER).  
Hänsyn tas till eventuella hål i polygonerna vid sammansmältningen.  
Denna operation är inte identisk med kombinera, som motsvarar en logisk XOR-operation.  
Dra ifrån  
Alla andra markerade polygoner dras bort från den polygon som ligger underst.  
Sedan subtraheras denna från den polygon som är placerad längst bak.  
Hänsyn tas till hål.  
Logiskt motsvarar den här operationen följande formel:  
A - (B1 _BAR_..... _BAR_ Bn)  
Skär av  
De markerade polygonerna sammanfattas till en enda polygon, som motsvarar snittmängden av alla ytor (logiskt OCH).  
Endast de ytor blir kvar där alla polygoner överlappar varandra.  
Visa diabild  
Här väljer du eller väljer bort en diabild för presentationen i diabildsvyn.  
Välj sedan menykommandot Bildskärmspresentation - Visa diabild eller klicka på ikonen Visa / dölj diabild på objektlisten.  
Du hittar även det här kommandot på den markerade diabildens snabbmeny.  
Diabildens rubrik (nere till höger om diabilden) får en grå bakgrund för att markera att denna diabild inte längre visas i presentationen.  
Genom att återigen välja menypunkten, eller genom att klicka på ikonen tar Du bort den grå bakgrunden och diabilden visas igen.  
Visa diabild  
Diabilder per rad  
Här anger du antalet diabilder per rad i diabildsvyn.  
Ju högre antal du väljer desto fler diabilder visas samtidigt på bildskärmen.  
Diabilder per rad  
Toningseffekt  
Toningseffekt  
Hastighet  
Hastighet  
Diabildsväxling  
Diabildsväxling  
Tid  
Tid  
Bildskärmspresentation med tidtagning  
Med det här kommandot startar du en presentation där visningstiden anges.  
Skillnaden jämfört med en "normal" presentation är att en klocka visas på bildskärmen.  
Under Presentationsinställningar... gör du standardinställningarna för en bildskärmspresentation.  
Bildskärmspresentation med tidtagning  
Aktuell storlek  
I detta fält på statuslisten finns information om markörens position och storleken på det aktuella objektet.  
Enheterna motsvarar enheterna på linjalerna.  
Du kan ställa in dem under Verktyg - Alternativ - Presentation - Allmänt.  
Aktuell sida / nivå  
I detta fält på statuslisten ser du det aktuella sidnumret i normalläget.  
Det visas i form av aktuellt sidnummer X och det total antalet sidor Y i dokumentet som Sida X / Y.  
Om Du har aktiverat nivåvyn ser Du här för varje aktiverat objekt på sidan namnet på nivån som innehåller objektet.  
Zoom  
Vid en lång klickning öppnar zoomningsverktyget fönstret Zooma.  
I det kan du ställa in vyskalan för bildskärmsvyn.  
Om du klickar kort aktiveras verktyget som visas i form av en ikon.  
Zoom  
Zoom (%PRODUCTNAME i dispositions - och diabildsvyn)  
Använd också tangentkombinationerna tangentkombinationerna tangentkombinationerna till att zooma.  
Förstora  
Detta verktyg används för att förstora vyn.  
Vyn förstoras med faktorn 2 när du klickar en gång.  
Istället för att klicka kan du också dra upp en rektangulär urvalsram.  
Ramens innehåll visas då formatfylld.  
Därefter kan verktyget inte längre aktiveras.  
Förstora  
Förminska  
Med detta verktyg förminskar Du vyn på bildskärmen med faktor 2.  
Därefter kan verktyget inte längre aktiveras.  
Förminska  
Zoom 100%  
Klicka på denna symbol för att ställa in vyn på bildskärmen på real storlek.  
Det innebär att 1 cm på bildskärmen motsvarar ca 1 cm på pappersutskriften (beror bl a på bildskärmens storlek).  
Zoom 100%  
Förra bilden  
Om Du tidigare ändrat dokumentets zoomvy återgår Du med denna ikon till den senaste visningen.  
Klicka en gång på den för att ställa in den senast inställda vyskalan.  
Du kan också trycka på Kommando Ctrl +kommatecken.  
Förra bilden  
Nästa bild  
Om Du tidigare ändrat dokumentets zoomvyer och återgått till den tidigare visningen, återgår Du med denna ikon till nästa visning.  
Klicka en gång på den för att ställa in den senast inställda vyskalan.  
Du kan också trycka på Kommando Ctrl +punkt.  
Nästa bild  
Hela sidan  
Klicka på denna symbol för att se hela sidans vy.  
Vyn väljs på ett sådant sätt att hela sidan visas.  
Hela sidan  
Sidbredd  
Klicka på denna symbol för att se hela sidbreddens vy.  
Sidbredd  
Optimal  
Med denna symbol ställer Du in vyn på ett sådant sätt att alla objekt på den visade sidan i dokumentet visas med maximal storlek.  
Optimal  
Objektzoom  
Klicka här om Du vill se det / de markerade objekten i maximal storlek.  
Objektzoom  
Flytta  
Med denna ikon blir markören till en hand, med vilken Du kan förskjuta fönstrets innehåll.  
Om Du nu pekar på dokumentet, håller musknappen nedtryckt och sedan drar musen följer dokumentet handen, som om Du flyttar en bit papper.  
Så snart Du släpper musknappen är det senast använda verktyget tillgängligt.  
Flytta  
Effekt  
Ikonen på verktygslisten i %PRODUCTNAME Draw öppnar fönstret Effekter.  
Här redigerar du objekt med olika effekter.  
Effekter  
Markera ett eller flera objekt.  
Nu visas de underordnade ikonerna till ikonen Effekt.  
Håll ner musknappen, för muspekaren till en av ikonerna och släpp upp musknappen.  
Då blir ikonen aktuellt effektverktyg och ersätter den tidigare ikonen Effekt på ritverktygslisten.  
Du kan även släppa upp musknappen och sedan dra i fönstrets titellist tills en fönsterkontur följer med muspekaren.  
Släpp upp musknappen nu så visas det fritt flyttbara fönstret Effekter.  
Effektfönstret ligger kvar på bildskärmen tills Du stänger det med stängningsknappen.  
Rotera  
Då kan du föra muspekaren till ett av objektets handtag.  
Över de fyra handtagen i hörnorna blir den till en öppen cirkelbåge och över de fyra handtagen i mitten av sidorna blir den till en förvrängningsmarkör.  
I mitten av objektet visas rotationspunkten som du kan flytta med musen.  
Rotationen sker runt den här punkten.  
Det kan bara finnas en rotationspunkt åt gången per sida på din teckning eller presentation.  
Fördelen med det är att Du kan vrida flera objekt (även objekt som infogats i efterhand) runt den gemensamma rotationspunkten.  
Om Du dubbelklickar på ett objekt placeras bl.a. rotationspunkten i mitten av objektet.  
Rotera objektet på samma nivå som sidan genom att placera markören på ett av de fyra hörnen och sedan dra.  
Rotera i tredje dimensionen, vinkelrätt mot sidan, genom att placera markören på ett av handtagen i mitten av de fyra sidorna och dra.  
Vid 3D-rotation blir den punkt som är längst bort från handtaget på den motstående sidan tillfälligt till rotationspunkt.  
Rotera  
Spegelvänd  
Välj det här verktyget för att spegelvända det markerade objektet.  
Du ser spegellinjen med punkter i varje ände.  
Du kan flytta de här punkterna en och en till en annan plats och flytta hela linjen utan att riktningen ändras genom att dra i spegellinjen mellan punkterna.  
Objektet spegelvänds över spegellinjen när du drar en av objektets handtag över spegellinjen och släpper det.  
Spegelvänd  
Till 3D-rotationsobjekt  
Med det här verktyget kan Du omvandla ett 2D-objekt till ett 3D-rotationsobjekt.  
Om Du har markerat ett 2D-objekt kan Du vrida det kring rotationsaxeln så att ett 3D-rotationsobjekt bildas.  
Rita ett 2D-objekt, t ex en bézierkurva som utgör halva konturen för en schackpjäs.  
Klicka på Till 3D-rotationsobjekt.  
Nu visas en symmetriaxel som Du kan flytta med musen.  
I ändarna på symmetriaxeln fins det små cirklar, som Du kan flytta med musen så att axelns vinkel ändras.  
Flytta nu axeln ett stycke tills en streckad spegelbild av 2D-objektet syns på andra sidan.  
Nu bildas ett 3D-objekt.  
Om de överlappar varandra skapas inte något 3D-objekt.  
Till 3D-rotationsobjekt  
Sätt på cirkel (perspektiviskt)  
Med det här verktyget placerar du det markerade objektet i perspektiv på en cirkel.  
Markera objektet, klicka på det här verktyget och placera sedan markören på ett av objektets åtta handtag.  
Muspekaren visas som ett slags krona.  
När du släpper upp musknappen passas objektet in i den nya ramkonturen.  
Sätt på cirkel (perspektiv)  
Sätt på cirkel (snedställ)  
Med det här verktyget kan Du placera det markerade objektet snedställt längs en cirkel.  
Funktionen motsvarar den med perspektiv enligt ovan.  
Sätt på cirkel (snedställ)  
Förvräng  
Med det här verktyget kan Du förvränga det markerade objektet.  
Du kan endast förvränga polygoner eller bézierkurvor.  
Om objektet, som Du vill förvränga, inte är en polygon eller bézierkurva, frågar %PRODUCTNAME om Du vill omvandla objektet.  
Vid förvrängning, till skillnad mot snedställning, kan Du ändra objektets kantlängd.  
Förvräng  
Transparens  
Med det här verktyget kan du definiera en transparensgradient interaktivt.  
Transparensgradienten fungerar som en linjär färggradient med gråskalor, där svart motsvarar 0% transparens och vitt motsvarar 100% transparens.  
Alla färger, som du t.ex. att drar och släpper från färglisten, omvandlas automatiskt till gråskalor som bestämmer transparensgraden.  
Klicka utanför det markerade området för att tillämpa gradienten och avsluta det här läget.  
Använd Ångra-funktionen om du inte vill tillämpa gradienten.  
Info:  
Effekten Transparens visas inte förrän du placerar en bakgrund eller ett objekt bakom det transparenta objektet.  
Transparens  
Färggradient  
Med det här verktyget kan Du ändra färggradienten interaktivt hos ett markerat objekt som redan har en färggradient.  
Den befintliga färggradienten (se Format - Yta - Färggradienter) är gränssättande för på vilket sätt Du kan göra ändringar interaktivt.  
Beroende på typen av färggradient kan Du redigera vektorn och färgobjekten.  
Du kan t ex dra färger från färglisten och släppa dem på färgobjekten.  
Klicka utanför det markerade området för att tillämpa gradienten och avsluta det här läget.  
Använd Ångra-funktionen om Du inte vill tillämpa gradienten.  
Efter det att Du har valt det här verktyget visas två färgobjekt, som förbinds med en vektor, i det markerade objektet.  
Beroende på typen av färggradient kan Du flytta det ena eller båda färgobjekten.  
Du kan ändra färgen hos färgobjekten var för sig genom att dra en färg från färglisten (meny Visa - Symbollister - Färglist) till ett av färgobjekten.  
Färggradient  
Objektlisten Redigera fästpunkter  
Denna objektlist syns bara när Du har klickat på ikonen Redigera fästpunkter på alternativlisten.  
Fästpunkter är punkter som Du själv har definierat till vilka förbindelse fästs.  
Dessutom finns det alltid de fyra fördefinierade fästpunkterna i mitten på den omgivande rektangeln på sidan.  
Infoga punkt  
Klicka på ikonen om Du vill infoga fästpunkter.  
Därefter infogar Du en fästpunkt varje gång Du klickar i det markerade objektet i dokumentet.  
Om Du vill sluta infoga punkter klickar Du på ikonen igen.  
Infoga punkt  
Vänster  
När Du klickar på den här ikonen så kommer riktningen för den förbindelse som fästs här att vara från objektet och ut åt vänster.  
Detta gäller den aktuella fästpunkten.  
Då väljer %PRODUCTNAME Impress den bästa vägen för förbindelsen.  
Vänster  
Överst  
Klicka på den här ikonen om Du vill att riktningen för den förbindelse som fästs vid den aktuella fästpunkten ska vara från objektet och uppåt.  
Överst  
Höger  
Klicka på den här ikonen om Du vill att riktningen för den förbindelse som fästs vid den aktuella fästpunkten ska vara från objektet och åt höger.  
Höger  
Underst  
Klicka på den här ikonen om Du vill att riktningen för den förbindelse som fästs vid den aktuella fästpunkten ska vara från objektet och nedåt.  
Underst  
Anpassa position till objekt  
När Du ändrar dimensionerna för ett objekt med fästpunkter påverkar detta även fästpunkterna, om Du har aktiverat den här ikonen.  
Inaktivera ikonen om Du inte vill att den aktuella fästpunkten ska ändra sitt läge i förhållande till objektsidan, när Du ändrar objektets storlek.  
Då kan Du välja någon av följande ikoner för att bestämma i förhållande till vilken sida som den aktuella fästpunktens position inte ska ändras.  
Anpassa position till objekt  
Fixerad horisontellt till vänster  
Den aktuella fästpunktens avstånd till objektets vänsterkant kommer att vara samma som tidigare, när Du ändrar objektets storlek.  
Fixerad horisontellt till vänster  
Fixerad horisontellt centrerad  
Den aktuella fästpunkten kommer att vara horisontellt centrerad mellan objektkanterna, när Du har ändrat objektets storlek.  
Fixerad horisontellt centrerad  
Fixerad horisontellt till höger  
Den aktuella fästpunktens avstånd till objektets högerkant kommer att vara samma som tidigare, när Du ändrar objektets storlek.  
Fixerad horisontellt till höger  
Fixerad vertikalt överkant  
Den aktuella fästpunktens avstånd till objektets överkant kommer att vara samma som tidigare, när Du ändrar objektets storlek.  
Fixerad vertikalt överkant  
Fixerad vertikalt centrerad  
Den aktuella fästpunkten kommer att vara vertikalt centrerad mellan objektkanterna, när Du har ändrat objektets storlek.  
Fixerad vertikalt centrerad  
Fixerad vertikalt nederkant  
Den aktuella fästpunktens avstånd till objektets underkant kommer att vara samma som tidigare, när Du ändrar objektets storlek.  
Fixerad vertikalt nederkant  
Text  
Ikonen öppnar utrullningslisten Text.  
Här kan du integrera texter i dina grafiska objekt.  
Texterna står antingen i en egen ram, är kopplade med ett annat objekt eller ram eller så bildar de en förklaring.  
Text  
Med denna ikon infogar du en text på sidan.  
Klicka på ikonen och rita upp en ram med musen för texten i dokumentet.  
Ramhöjden är automatiskt enradig.  
Klicka på ikonen och rita upp en ram, som kommer att avgränsa texten, i dokumentet med musen.  
Runt om textramen ritas en skrafferad ram med vilken textobjektet kan förskjutas.  
Så snart du släpper musknappen är textmarkören klar för inmatning av texten.  
Klicka utanför textramen för att avsluta textinmatningen.  
Du kan senare redigera texten genom att helt enkelt klicka på den.  
Text  
Anpassa text till ram  
Den här ikonen används för att mata in en text, vars teckenstorlek är kopplad till ramens storlek.  
Klicka på ikonen och rita upp en ram som avgränsar texten i dokumentet med musen.  
Mata nu in texten.  
Klicka utanför textramen för att avsluta textinmatningen.  
Du kan redigera texten senare genom att helt enkelt klicka på den.  
Om ramen flyttas, kopieras eller raderas, gäller det också den kopplade texten.  
Anpassa text till ram  
Förklaring  
Med denna ikon skriver Du in en förklaring.  
Klicka först på ikonen och sedan på det ställe i dokumentet som pekaren ska peka på.  
Håll musknappen nedtryckt och dra till det ställe där förklaringstexten ska visas.  
Släpp musknappen.  
Klicka sedan i textfältet.  
Mata nu in texten.  
Fältet med förklaringstexten förstoras automatiskt upp till en viss storlek om Du matar in mer text.  
Om texten inte ryms i den förinmatade storleken radbryts den med hänsyn till avstavningsreglerna.  
Generellt sett försöker programmet göra en radbrytning utan att dela orden.  
Förklaring  
Om Du i redigeringsläget klickar på textens grå ram, lämnar Du läget.  
Om Du vill, kan Du omedelbart radera objektet med tangenten Delete.  
Anpassa vertikal text till ram  
Med den här ikonen kan du skriva en vertikal text vars teckenstorlek är kopplad till storleken på textens ram  
Anpassa vertikal text till ram  
Rektanglar  
Utrullningslisten Rektanglar innehåller fyllda och tomma former som du kan infoga på sidan.  
Klicka på önskad symbol och dra upp en rektangel på sidan.  
Den fylls med önskat innehåll.  
Via menyn Format eller snabbmenyn kan du sedan använda kommandona för formatering och ändring av objektet.  
Rektangel  
Med den här funktionen ritar du en fylld rektangel.  
Rektangel  
Kvadrat  
Här ritar du upp en fylld kvadrat.  
Kvadrat  
Rundad rektangel  
Med den här funktionen ritar Du en rundad, fylld rektangel.  
Rundad rektangel  
Rundad kvadrat  
Med den här funktionen ritar Du en rundad, fylld kvadrat.  
Rundad kvadrat  
Ofylld rektangel  
Med den här funktionen ritar Du en ofylld rektangel.  
Rektangel, ofylld  
Ofylld kvadrat  
Med den här funktionen ritar Du en ofylld kvadrat.  
Kvadrat, ofylld  
Rundad rektangel, ofylld  
Med den här funktionen ritar Du en rundad, ofylld rektangel.  
Rundad rektangel, ofylld  
Rundad kvadrat, ofylld  
Med den här funktionen ritar Du en rundad, ofylld kvadrat.  
Rundad kvadrat, ofylld  
Ellipser  
Utrullningslisten Ellipser innehåller ellipser och cirklar som du kan infoga på sidan.  
Klicka på önskad symbol och dra upp en rektangel på sidan.  
Den fylls med önskat innehåll.  
Rita först en cirkel eller ellips och släpp därefter musknappen.  
Nu visas en radie i objektet som följer varje musrörelse.  
Klicka en gång när radien motsvarar radien för önskad sektor, segment eller båge.  
En ny radie följer musens rörelse.  
Klicka åter en gång när radien motsvarar den andra radien.  
Du kan också begränsa radiens vinkel till 45 grader.  
Ellips  
Här ritar du upp en fylld ellips genom att dra med musen.  
Ellips  
Cirkel  
Här ritar du upp en fylld cirkel genom att dra med musen.  
Cirkel  
Ellipssektor  
Här ritar du upp en fylld ellipssektor genom att dra med musen.  
Ellipssektor  
Cirkelsektor  
Här ritar du upp en fylld cirkelsektor genom att dra med musen.  
Cirkelsektor  
Ellipssegment  
Här ritar du upp ett fyllt ellipssegment genom att dra med musen.  
Ellipssegment  
Cirkelsegment  
Här ritar du upp ett fyllt cirkelsegment genom att dra med musen.  
Cirkelsegment  
Ellips, ofylld  
Här ritar du upp en ofylld ellips genom att dra med musen.  
Ellips, ofylld  
Cirkel, ofylld  
Här ritar du upp en ofylld cirkel genom att dra med musen.  
Cirkel, ofylld  
Ellipssektor, ofylld  
Här ritar du upp en ofylld ellipssektor genom att dra med musen.  
Ellipssektor, ofylld  
Cirkelsektor, ofylld  
Här ritar du upp en ofylld cirkelsektor genom att dra med musen.  
Cirkelsektor, ofylld  
Ellipssegment, ofyllt  
Här ritar du upp ett ofyllt ellipssegment genom att dra med musen.  
Ellipssegment, ofyllt  
Cirkelsegment, ofyllt  
Här ritar du upp ett ofyllt cirkelsegment genom att dra med musen.  
Cirkelsegment, ofyllt  
Ellipsbåge  
Här ritar du upp en ellipsbåge genom att dra med musen.  
Ellipsbåge  
Cirkelbåge  
Här ritar du upp en cirkelbåge.  
Cirkelbåge  
Kurvor  
Utrullningslisten Kurvor innehåller ikoner som används till att rita kurvor.  
Genom att hålla skifttangenten nedtryckt begränsar Du musens rörelse till multiplar av 45 grader.  
Då kan Du skapa objekt som kombineras av kurvor som inte hänger ihop.  
Det blir alltså ett hål i det större objektet.  
Kurva, fylld  
Klicka på ikonen.  
Nu kan du definiera en kurva i dokumentet genom att definiera tre stödpunkter.  
Kurvan kommer att följa musens rörelse så gott det går.  
Definiera stödpunkter genom att klicka med musen och bestäm andra delar av kurvan genom att dra med musen.  
Kurvan fylls automatiskt med den aktuella ytfärgen.  
Via kurvans snabbmeny kan Du förstås välja att i stället fylla den med en färggradient, en bitmap eller en skraffering.  
Kurva, fylld  
Polygon, fylld  
Klicka på ikonen.  
Definiera nu polygonens punkter genom att först rita upp en linje i dokumentet för att fastlägga de första två punkterna.  
De andra punkterna definierar Du genom att klicka i dokumentet.  
Punkterna förbinds med räta linjer.  
Genom att dubbelklicka sluter Du polygonen som fylls automatiskt.  
Polygon, fylld  
Polygon (45°), fylld  
Med denna ikon ritar Du en fylld polygon.  
Vinklarna är begränsade till multiplar av 45 grader, med undantag av den sista linjen som sluter polygonen.  
Klicka på ikonen.  
Definiera nu polygonens punkter genom att först rita upp en linje i dokumentet för att fastlägga de första två punkterna.  
De andra punkterna definierar Du genom att klicka i dokumentet.  
Punkterna förbinds med räta linjer.  
Genom att dubbelklicka sluter Du polygonen som fylls automatiskt.  
Polygon (45°), fylld  
Frihandslinje  
Med den här ikonen definierar Du en fylld, frihandslinje.  
Rita nu en valfri linje med musknappen nedtryckt.  
När Du släpper musknappen sluts linjen automatiskt med hjälp av en rät linje som %PRODUCTNAME automatiskt skapar.  
Ytan mellan linjerna fylls med den aktuella ytfärgen.  
Frihandslinje  
Kurva  
Kurva  
Klicka på ikonen.  
Nu kan Du definiera en kurva på sidan genom att klicka på tre stödpunkter.  
När Du klickar på den tredje punkten beräknar programmet bézierkurvan och visar den.  
Polygon  
Polygon  
Polygon (45°)  
Med denna ikon ritar Du en polygon.  
Vinklarna är begränsade till multiplar av 45 grader, med undantag av den sista linjen som sluter polygonen.  
Definiera nu polygonpunkterna genom att klicka på sidan.  
Punkterna förbinds med räta linjer.  
Du kan också infoga valfria delar av polygonen genom att dra med musen.  
Dessa sätts då in i 45 graders vinkel som korta linjer.  
Däremot fylls den inte.  
Polygon (45°)  
Frihandskurva  
Frihandskurva  
3D-objekt  
Utrullningslisten 3D-objekt använder du när du vill rita 3D-objekt.  
Dra sedan upp en ram i önskad objektstorlek på sidan.  
Så snart du släpper musknappen ritas 3D-objektet.  
3D-objekt öppnas alltid med lika långa sidor, alltså t.ex. som kub eller klot.  
Om du inte vill det kan du hålla ner skifttangenten när du först ritar upp ett 3D-objekt.  
3D-objekt  
3D-objekt kan placeras och roteras valfritt i rummet.  
För att rotera använder du rotationsverktyget på utrullningslisten Effekter.  
Kub  
Med den här ikonen definierar du en 3D-kub.  
Kub  
Klot  
Den här ikonen definierar ett klot.  
Klotet har två poler, som är förbundna med längdgraderna och ett antal breddgrader.  
Du ser den här indelningen om du växlar linjestilen i listrutan med samma namn till t.ex. "Genomgående".  
Klot  
Cylinder  
Med den här ikonen infogar du en cylinder.  
Cylinder  
Kon  
Med den här ikonen infogar du en kon.  
Kon  
Pyramid  
Med denna ikon infogar du en pyramid med fyra grundkanter.  
Om du t.ex. vill ha en pyramid med en trekantig bottenyta kan du ange 3 i fönstret 3D-effekter - Geometri - Segment - Horisontell.  
Pyramid  
Torus  
Med den här ikonen infogar du en torus.  
Torus  
Skal  
Med den här ikonen infogar du ett skal.  
Skal  
Halvklot  
Med den här ikonen infogar du ett halvklot.  
Halvklot  
Förbindelse  
Förbindelse används till att koppla ihop objekt med en linje.  
Om du flyttar objekten anpassas förbindelsen automatiskt.  
Vid kopiering av ihopkopplade objekt kopieras även förbindelserna.  
Förbindelse  
Klicka på ikonen.  
Muspekaren får nu förbindelsens tecken, ända tills Du avslutar förbindelseläget.  
Du kan nu koppla samman två objekt med en linje genom att dra musen från det ena till det andra objektet.  
Om Du i efterhand vid ändra Förbindelsens egenskaper har Du diverse olika möjligheter att göra detta under Format.  
I annat fall måste Du sätta musen på kanten av objektet.  
Du ser nu att objektet blinkar med regelbundna intervall.  
Håll musknappen nedtryckt och drag till det andra objektet.  
Även här pekar Du antingen mitt i eller på kanten, tills objektet börjar blinka.  
Båda objekt är nu förbundna med varandra.  
Vid den beskrivna metoden letar %PRODUCTNAME själv rätt på den optimala punkten för att fästa förbindelsen under den omgivande rektangelns fyra sidors mittpunkter.  
Om du själv vill bestämma den sida vid vilken förbindelsen ska fästas, för du muspekaren till exakt mitten av den omgivande rektangelns aktuella sida.  
Här börjar nu en liten kvadrat att blinka.  
Denna metod, med vilken Du fäster förbindelsen på mitten av en av den omgivande rektangelns sidor, är dock bara användbar för rektangulära objekt.  
Vid ellipser eller oregelbundna objekt blir förbindelsen för det mesta felplacerad på den omgivande rektangeln.  
Inom den omgivande rektangeln kan Du definiera godtyckliga fästpunkter vid vilka förbindelserna kan fästas med fästpunktsredigeraren, som Du hittar på utrullningslisten, Effekter.  
Du kan redigera förbindelserna (t ex linjestil, linjeslut och färger) - se Objektlist) och radera (markera och tryck tangenten Delete).  
Förbindelse  
Med denna ikon infogar Du en förbindelse.  
Förbindelse  
Förbindelsen börjar med en pilspets  
Med denna ikon infogar Du en förbindelse som börjar med en pilspets.  
Förbindelsen börjar med en pilspets  
Förbindelsen slutar med en pilspets  
Med denna ikon infogar Du en förbindelse som slutar med en pilspets.  
Förbindelsen slutar med en pilspets  
Förbindelse med pilspetsar  
Med denna ikon infogar Du en förbindelse med pilspetsar.  
Förbindelse med pilspetsar  
Förbindelsen börjar med en cirkel  
Med denna ikon infogar Du en förbindelse som börjar med en cirkel.  
Förbindelsen börjar med en cirkel  
Förbindelse slutar med cirkel  
Med denna ikon infogar Du en förbindelse som slutar med en cirkel.  
Förbindelsen slutar med en cirkel  
Förbindelse med cirklar  
Med denna ikon infogar Du en förbindelse med cirklar.  
Förbindelse med cirklar  
Förbindelselinje  
Med denna ikon infogar Du en förbindelselinje.  
Förbindelselinje  
Förbindelselinjen börjar med en pilspets  
Med denna ikon infogar Du en förbindelselinje som börjar med en pilspets.  
Förbindelselinjen börjar med en pilspets  
Förbindelselinje slutar med pilspets  
Med denna ikon infogar Du en förbindelselinje som slutar med en pilspets.  
Förbindelselinjen slutar med en pilspets  
Förbindelselinje med pilspetsar  
Med denna ikon infogar Du en förbindelselinje med pilspetsar.  
Förbindelselinje med pilspetsar  
Förbindelselinjen börjar med en cirkel  
Med denna ikon infogar Du en förbindelselinje som börjar med en cirkel.  
Förbindelselinje börjar med cirkel  
Förbindelselinjen slutar med en cirkel  
Med denna ikon infogar Du en förbindelselinje som slutar med en cirkel.  
Förbindelselinjen slutar med en cirkel  
Förbindelselinje med cirklar  
Med denna ikon infogar Du en förbindelselinje med cirklar.  
Förbindelselinje med cirklar  
Direktförbindelse  
Med denna ikon infogar Du en direktförbindelse.  
Direktförbindelse  
Direktförbindelsen börjar med en pilspets  
Med denna ikon infogar Du en direktförbindelse som börjar med en pilspets.  
Direktförbindelsen börjar med en pilspets  
Direktförbindelsen slutar med en pilspets  
Med denna ikon infogar Du en direktförbindelse som slutar med en pilspets.  
Direktförbindelsen slutar med en pilspets  
Direktförbindelse med pilspetsar  
Med denna ikon infogar Du en direktförbindelse med pilspetsar.  
Direktförbindelse med pilspetsar  
Direktförbindelsen börjar med en cirkel  
Med denna ikon infogar Du en direktförbindelse som börjar med en cirkel.  
Direktförbindelsen börjar med en cirkel  
Direktförbindelsen slutar med en cirkel  
Med denna ikon infogar Du en direktförbindelse som slutar med en cirkel.  
Direktförbindelsen slutar med en cirkel  
Direktförbindelse med cirklar  
Med denna ikon infogar Du en direktförbindelse med cirklar.  
Direktförbindelse med cirklar  
Kurvförbindelse  
Med denna ikon infogar Du en kurvförbindelse.  
Kurvförbindelse  
Kurvförbindelsen börjar med en pilspets  
Med denna ikon infogar Du en direktförbindelse med pilspets.  
Kurvförbindelsen börjar med en pilspets  
Kurvförbindelse slutar med pilspets  
Med denna ikon infogar Du en kurvförbindelse som slutar med en pilspets.  
Kurvförbindelsen slutar med en pilspets  
Kurvförbindelse med pilspetsar  
Med denna ikon infogar Du en kurvförbindelse med pilspetsar.  
Kurvförbindelse med pilspetsar  
Kurvförbindelsen börjar med en cirkel  
Med denna ikon infogar Du en kurvförbindelse som börjar med en cirkel.  
Kurvförbindelse börjar med cirkel  
Kurvförbindelse slutar med cirkel  
Med denna ikon infogar Du en kurvförbindelse som slutar med en cirkel.  
Kurvförbindelsen slutar med en cirkel  
Kurvförbindelse med cirklar  
Med denna ikon infogar Du en kurvförbindelse med cirklar.  
Kurvförbindelse med cirklar  
Infoga  
Med den här ikonen öppnar du en utrullningslist med funktioner för att infoga diagram, grafikobjekt, tabeller, filer, bilder och sidor.  
Ikon på verktygslisten:  
Infoga  
När Du en gång har valt en funktion på utrullningslisten, visas alltid ikonen för den senast infogade funktionen.  
Du kan nu upprepa den senast funktionen genom att klicka snabbt, eller öppna utrullningslisten igen genom att klicka litet längre.  
Infoga diagram  
Infoga formel  
Infoga ram  
Infoga OLE-objekt  
Infoga PlugIn  
Infoga Applet  
Infoga %PRODUCTNAME Calc-tabell  
Fil  
Infoga sida  
Infoga grafik  
Infoga ljud-PlugIn  
Infoga video-PlugIn  
Linjer och pilar  
Utrullningslisten Linjer och pilar innehåller ikoner som används till att rita linjer med olika slut.  
Linjesluten kan du också definiera senare.  
I så fall väljer du kommandot Linje på t.ex. snabbmenyn till den / de markerade linjen / linjerna.  
Linjer och pilar  
Linje  
Med denna ikon ritar Du en rak linje utan framhävda linjeslut.  
Linje  
Linje med pilslut  
Med denna ikon ritar Du en rak linje som slutar med en pilspets.  
Linje med pilslut  
Linje med pil - / cirkelslut  
Med denna ikon ritar Du en rak linje som börjar med en pilspets och slutar med en cirkel.  
Linje med pil - / cirkelslut  
Linje med pil - / kvadratslut  
Med denna ikon ritar Du en rak linje som börjar med en pilspets och slutar med en kvadrat.  
Linje med pil - / kvadratslut  
Linje (45°)  
Med denna ikon ritar Du en rak linje med en vinkel på 45 grader.  
Linje (45°)  
Linje med pilbörjan  
Med denna ikon ritar Du en rak linje som börjar med en pilspets.  
Linje med pilbörjan  
Linje med cirkel - / pilslut  
Med denna ikon ritar Du en rak linje som börjar med en cirkel och slutar med en pilspets.  
Linje med cirkel - / pilslut  
Linje med kvadrat - / pilslut  
Med denna ikon ritar Du en rak linje som börjar med en kvadrat och slutar med en pilspets.  
Linje med kvadrat - / pilslut  
Måttlinje  
Med denna ikon drar Du upp en måttlinje Klicka på ikonen.  
Definiera ny begynnelsepunkt för Din dimensioneringslinje genom att trycka med musknappen där.  
Håll musknappen nedtryckt och dra upp måttlinjen.  
Släpp musknappen där måttlinjen ska sluta.  
Håll ner skifttangenten när Du drar upp måttlinjen för att göra måttlinjen exakt horisontell eller vertikal eller i 45 graders vinkel.  
Håll ner Kommando Ctrl -tangenten för att låta måttlinjen börja och sluta exakt vid de närmast liggande objektsidorna.  
Tänk dock på att måttsättningstalet vid storleksförändringar inte längre ändras automatiskt efter omvandling till polygoner, utan förblir detsamma.  
Ytterligare information finns i hjälpen till menykommandot Format - Dimensionering.  
Måttlinje  
Linje med pilslut  
Med denna ikon ritar Du en rak linje med som börjar och slutar med pilspetsar.  
Linje med pilslut  
3D-effekter  
Med ikonen 3D-controller visar du fönstret 3D-effekter där du skapar och redigerar 3D-objekt.  
Du kan skapa ett 3D-objekt av ett eller flera markerade 2D-objekt och sedan tilldela detta 3D-objekt egenskaper.  
Du kan t.ex. bestämma antal, position, färg och ljusstyrka hos ljuskällorna som lyser på 3D-objektet.  
Du kan låta det här fönstret vara öppet medan du redigerar dokumentet.  
Det är också åtkomligt via menykommandot Format - 3D-effekter.  
3D-controller  
Första nivån  
Med den här ikonen döljer du alla nivåer som står under den första nivån i hierarkin.  
Om du vill visa alla nivåer igen klickar du på ikonen Alla nivåer.  
Första nivån  
Alla nivåer  
Med denna ikon visar du alla nivåer som du tidigare dolt med kommandot Första nivån.  
Alla nivåer  
Dölj understycken  
Med den här ikonen döljer du alla element som finns under den aktuella nivån i hierarkin.  
Om du vill visa nivåerna igen klickar du på ikonen Visa understycken.  
Dölj understycken  
Visa understycken  
Med denna ikon visar du alla nivåer som du tidigare dolt med kommandot Dölj understycken.  
Visa understycken  
Formatering på / av  
Med den här ikonen växlar du textvyn i dispositionen mellan "formaterad" (med textattribut som på diabilden) och "oformaterad ".  
Du kan ändra standardinställningarna för formateringen i Stylist genom att där öppna snabbmenyn till en presentationsobjektmall och klicka på Ändra.  
Formatering på / av  
Svartvit-vy  
Med den här ikonen växlar Du mellan att visa texten i svartvitt eller i färg i dispositionsvyn.  
Antingen visas texterna i dispositionen bara i svartvitt eller så har de samma färg som på diabilden.  
Svartvit-vy  
Redigera fästpunkter  
Med det här verktyget kan du redigera fästpunkterna för ett markerat objekt.  
Till fästpunkterna kan du t.ex. ansluta förbindelser.  
När du har valt verktyget visas fler ikoner för redigering av fästpunkterna på objektlisten.  
Redigera fästpunkter  
Rotationsläge efter klick på objekt  
Med den här funktionen tilldelas ett objekt rotationsläge när du har klickat på det två gånger.  
Du kan rotera objektet i valfri vinkel genom att dra i ett av handtagen.  
Rotationsläge efter klick på objekt  
Tillåta effekter  
Om du aktiverar den här funktionen visas de tilldelade effekterna direkt i dokumentet utan att du behöver starta en presentation.  
Om du pekar med musen på ett objekt som tilldelats en effekt så ändrar muspekaren utseende till en hand med ett pekfinger.  
Om du klickar då så tillämpas effekten.  
Om du vill klicka på objektet för att redigera det måste du hålla ned Alternativ Alt -tangenten när du klickar.  
Tillåt effekter  
Tillåt interaktioner  
Om du aktiverar den här ikonen kan du utföra interaktioner direkt i dokumentet utan att behöva starta en presentation.  
Du kan tilldela ett objekt interaktioner via menyn Bildskärmspresentation - Interaktion....  
Du kan t.ex. hoppa till nästa sida, eller köra ett makro genom att klicka på ett grafikobjekt.  
Om du pekar med musen på ett objekt som tilldelats en interaktion så ändrar muspekaren utseende till en hand med ett pekfinger.  
Om du klickar då så utförs interaktionen.  
Om du vill klicka på objektet för att redigera det måste du hålla ned Alternativ Alt -tangenten när du klickar.  
Under en löpande presentation förblir dock objektet osynligt.  
Tillåt interaktion  
Visa stödlinjer  
Om du aktiverar den här ikonen visas stödlinjerna på bildskärmen.  
När ikonen inte är aktiverad är stödlinjerna osynliga men fungerar ändå.  
Visa stödlinjer  
Dubbelklicka för att redigera text  
Om du aktiverar den här ikonen kan du växla direkt till textredigeringsläget genom att dubbelklicka på ett textobjekt.  
Du kan då skriva över, ändra eller radera text.  
Dubbelklicka för att redigera text  
Enkla handtag  
Med den här ikonen kan du definiera att markerade objekt ska ha enkla 2D-handtag.  
Handtagen visas som plana ytor utan 3D-effekt.  
Enkla handtag  
Stora handtag  
Om du klickar på den här ikonen visas handtagen förstorade.  
Då blir det lättare att "ta tag" i handtagen med musen.  
Stora handtag  
Skapa objekt med attribut  
Om du klickar på den här ikonen fylls objekt med attribut när du ritar upp dem.  
Du kan t.ex. välja en färggradient och en inramningsfärg på objektlisten.  
Om du sedan ritar upp en rektangel fylls den direkt med de valda attributen.  
Skapa objekt med attribut  
Lämna alla grupperingar  
Klicka på den här ikonen om du vill lämna alla grupperingar.  
Den här ikonen är bara tillgänglig om du har gått in i en gruppering.  
Lämna alla grupperingar  
Fäst mot stödlinjer  
Fäst mot stödlinjer  
Fäst mot sidmarginaler  
Fäst mot sidmarginaler  
Fäst mot objektram  
Fäst mot objektram  
Fäst mot objektpunkter  
Fäst mot objektpunkter  
Tillåt snabbredigering  
Tillåt snabbredigering  
Bara textområde kan markeras  
Bara textområde kan markeras  
Antyd extern grafik  
Antyd extern grafik  
Konturläge  
Konturläge  
Antyd text  
Inga fyllningar  
Visa bara fina linjer  
Visa bara fina linjer  
Kortkommandon för presentationsdokument  
Här hittar du tangentkombinationer som du kan använda i presentationsdokument.  
Dessutom gäller de allmänna tangentkombinationerna i %PRODUCTNAME.  
Funktionstangenter vid presentationsdokument  
Tangentkombination  
Effekt  
F2  
Redigera text  
Kommando Ctrl +F2  
Bildskärmspresentation  
F3  
Gå in i gruppering  
Kommando Ctrl +F3  
Lämna gruppering  
Skift+F3  
Duplicera  
F4  
Position och storlek  
F5  
Navigator  
F7  
Rättstavningskontroll  
Kommando Ctrl +F7  
Synonymordlista  
F8  
Redigera punkter  
Kommando Ctrl +Skift+F8  
Anpassa text till ram  
F11  
Stylist  
F12  
Dispositionsvy  
Kommando Ctrl  
Teckningsvy  
Tangentstyrning vid presentationer  
Tangentkombination  
Effekt  
Esc  
Avsluta presentation  
Blankstegstangenten  
Nästa objektanimation resp. nästa diabild  
Returtangenten  
Nästa diabild  
nn returtangenten  
Växla diabild till den nn:te diabilden  
Vänsterpilstangenten  
Växla diabild till föregående diabild  
Högerpilstangenten  
Växla diabild till nästa diabild  
Home  
Växla diabild till första diabilden  
End  
Växla diabild till sista diabilden  
PageUp  
Växla till föregående sida  
PageDown  
Växla till nästa sida  
F5  
Öppna Navigator  
Tangentstyrning i teckningsvyn  
Tangentkombination  
Effekt  
PageUp  
Växla till föregående sida  
PageDown  
Växla till nästa sida  
+ tangent  
Förstorar vyn  
- tangent  
Förminskar vyn  
×-tangent (numeriska tangentbordet)  
Zoom till den aktuella markeringen  
÷-tangent (numeriska tangentbordet)  
Zoom på hela sidan  
Kommando Ctrl +G  
Gruppering / Gruppera  
Skift + Kommando+Alternativ Ctrl+Alt +A  
Upphäv gruppering  
Nedtryckt Skift - vänster musknapp  
Sammanställ gruppering, skifttangenten ska hållas ner tills markeringen av objekt med musklick har avslutats.  
Nedtryckt Kommando Ctrl - vänster mustangent  
Redigera gruppering, d.v.s. markera enskilda objekt i en gruppering genom att klicka med musen.  
Kommando Ctrl +K  
Kombination  
Skift + Kommando+Alternativ Ctrl+Alt +K  
Upphäv kombination  
Skift + Kommando Ctrl och +  
Längst fram  
Kommando Ctrl och +  
Längre fram  
Kommando Ctrl och -  
Längre bak  
Skift + Kommando Ctrl och -  
Längst bak  
Speciella tangentstyrningar vid presentationsdokument  
Tangentkombination  
Effekt  
Piltangent  
Flyttar det markerade objektet i pilens riktning.  
Kommando Ctrl och piltangent  
Flyttar sidvyn i önskad riktning.  
Nedtryckt skifttangent och dra med musen  
Det markerade objektet flyttas exakt horisontellt eller vertikalt i den önskade riktningen.  
Kommando Ctrl och dra med mus och aktivt alternativ Kopia vid flyttning  
När du flyttar det markerade objektet skapas en kopia.  
Alternativ Alt  
När objekt skapas eller när deras storlek ändras, centreras de efter att tangenten Alternativ Alt tryckts.  
Alternativ Alt och klicka med musen på objekt  
Markering av överlappande objekt.  
Objektet som ligger bakom det markerade objektet markeras.  
Alternativ Alt +Skift och klicka med musen på objekt  
Markering av överlappande objekt.  
Objektet som ligger framför det markerade objektet markeras.  
Skifttangent vid markering av objekt  
Objekt tillfogas markeringen om det ännu inte markerats, eller tas bort från markeringen om det redan varit markerat innan.  
Skifttangent vid förstora / skapa  
Objekt förstoras proportionellt mot ursprungsformen.  
En rak linje kan bara ändras i sin riktning.  
Tabbtangent  
Det görs en markering av de enskilda objekten i den ordning de skapats, från det första till det sista objektet.  
Skift+tabbtangent  
Markering av objekten i den ordning de skapades, från det sista till det första objektet.  
Skifttangent när musen dras i läget Redigera punkter  
Gör det möjligt att ändra en måttlinjes längd.  
Esc-tangent  
Skiftar till markeringsläget när ett skapa-verktyg är aktivt.  
Stänger av markeringen när ett objekt markerats.  
Skiftar tillbaka ett objekt, som står i textinmatningsläget, från textinmatningsläget.  
Objektet fortsätter att vara markerat  
Omvandla till kurva, polygon, 3D  
Många objekt kan du redigera mycket effektfullt med en omvandling.  
Prova själv!  
Här följer ett mycket enkelt exempel som visar vad du kan göra.  
Rita upp en rektangel med musen.  
Den har standardinställningarna för färg, linjetjocklek, o.s.v. och bör nu vara markerad.  
Välj Ändra - Omvandla. (I %PRODUCTNAME Impress hittar du motsvarande kommando på snabbmenyn till rektangeln.) Du ser bl.a. följande kommandon på undermenyn:  
Till kurva, Till polygon, Till 3D, Till 3D-rotationsobjekt.  
Med kommandot Ändra - Omvandla - Till kurva omvandlar du rektangeln till en Bézierkurva.  
Nu kan du redigera punkterna.  
Du kan flytta dem, omvandla dem från hörnpunkt till rundad punkt, radera dem, infoga nya punkter och så vidare.  
Alla möjligheter beskrivs utförligt till sökorden Punkter, redigera och Bézierobjektlist i %PRODUCTNAME -hjälpen.  
Med kommandot Ändra - Omvandla - Till polygon omvandlar du den ursprungliga rektangeln till en "polygon med 4 punkter" vilket du kan läsa efteråt i statuslisten.  
Du kan nu t.ex. bryta ner polygonen till sina grundläggande beståndsdelar.  
Kommandot finns på menyn Ändra och heter Bryt ner.  
Statuslisten visar sedan "4 linjer".  
De här linjerna kan du flytta på en och en.  
Dessutom kan du också markera polygonen och ändra punkter, infoga nya o.s.v. med ikonen Redigera punkter.  
Med kommandot Ändra - Omvandla - Till 3D skapar du ett tredimensionellt objekt av ett tvådimensionellt objekt med en såkallad extrusion.  
Polygonen "dras" lodrätt i förhållande till sin yta till den tredje dimensionen.  
3D-objektet kan du rotera fritt och redigera med hjälp av fönstret 3D-effekter som du kan öppna från snabbmenyn.  
Med kommandot Ändra - Omvandla - Till 3D-rotationsobjekt skapar du ett 3D-objekt med en såkallad roteringsextrusion.  
En polygon roteras med 360 grader runt en axel till den tredje dimensionen.  
Om du roterar rektangeln något innan den omvandlas till ett 3D-rotationsobjekt, skapar du ett ännu mer iögonfallande objekt.  
Skapa animerad GIF-bild  
Du kan även skapa rörliga bilder, d.v.s. små tecknade filmer, till dina presentationer och spela upp dem.  
Du kan använda animationsformatet i %PRODUCTNAME Impress.  
Dessutom kan du visa animerade GIF-bilder.  
Du kan dra dem till dina dokument med musen.  
Animerade GIF-bilder är ett utmärkt sätt att väcka intresse för Internetsidor och andra presentationer.  
En animerad GIF-bild består av en serie av pixelbilder som på ett mycket utrymmessnålt sätt har placerats i en enda fil.  
Dessa laddas till arbetsminnet och kan sedan visas av något program som kan hantera animerade GIF-bilder, t.ex. de flesta webbläsare och givetvis även %PRODUCTNAME.  
Om du väljer att visa den animerade GIF-bilden så att flera bilder per sekund upprepas i en ändlös slinga, uppfattas bilderna som små tecknade filmer.  
Innan du kan sammanställa en animation, måste du först rita alla enskilda bilder.  
I det här exemplet används en toning för att du inte ska behöva rita alla de enskilda bilderna.  
I följande exempel används en toning för att du snabbt ska få ihop tio eller fler enstaka bilder till animationen.  
Eftersom en toning bara kan utföras i %PRODUCTNAME Draw, en animation däremot bara i %PRODUCTNAME Impress, används ett teckningsdokument och ett presentationsdokument i det här exemplet.  
Öppna ett nytt tomt teckningsdokument (Nytt - Teckning).  
Rita t.ex. en röd fylld rektangel uppe till vänster och en grön fylld cirkel nere till höger.  
Markera båda objekten (håll ner skifttangenten).  
Välj Redigera - Tona över.  
I dialogrutan väljer du 8 steg och Tona över attribut.  
Klicka på OK.  
Du ser nu 10 objekt som bildar en grupp.  
I så fall behåller du grupperingen.  
Om du däremot vill att den animerade GIF-bilden ska visa ett centrerat objekt som fyller hela bilden och ändrar sin form och färg, men inte förflyttar sig uppe från vänster ner till höger tvärs över bilden, ska du nu upphäva grupperingen (i menyn Ändra).  
I det här exemplet har grupperingen upphävts (Ändra - Upphäv gruppering).  
Kopiera nu alla enstaka bilder tillsammans (de är fortfarande gemensamt markerade) till urklippet.  
Växla till ett tomt presentationsdokument i %PRODUCTNAME Impress.  
Där klistrar du in innehållet från urklippet.  
Nu ska du fortsätta arbetet i %PRODUCTNAME Impress, eftersom alla enskilda bilder har skapats.  
Välj kommandot Bildskärmspresentation - Animation.  
Dialogrutan Animation visas.  
Välj alternativet Bitmapobjekt.  
GIF-bilder är bitmap - eller pixelbilder.  
Alla enskilda objekt är fortfarande markerade (och ligger i rätt ordning ovanpå varandra).  
Klicka på ikonen Överta objekt ett och ett.  
De 10 enskilda objekten överförs som bitmaps i 10 bilder i animationen.  
Objektet längst bak eller längst ned i stapeln används till bild 1, det översta till bild 10.  
Du kan titta på resultatet i dialogrutan (symbolen Spela upp).  
Om animationen ska spelas upp med bra flyt, är det vara bättre att den spelar bild 10, via 9, 8 och så vidare tillbaka till bild 2.  
Sedan visas hela bildserien igen, med start från bild 1.  
Gör så här:  
1.  
Se till att bild 10 i dialogrutan Animation är aktuell bild (ikonen Sista bilden).  
Markera som enda objekt det näst sista objektet före den gröna cirkeln ("objekt från bild 9") i presentationsdokumentet (du ska inte ändra något i dialogrutan Animation!).  
Klicka sedan på ikonen Överta objekt i dialogrutan Animation.  
2.  
Markera nästa objekt ("objekt till bild 8"), och klicka på Överta objekt i dialogrutan Animation.  
Fortsätt sedan på samma sätt ända fram till "objekt till Bild 2", det andra objektet uppe till vänster.  
3.  
Nu kan du överföra den färdiga animationen till sidan genom att klicka på kommandoknappen Skapa.  
4.  
Det animerade bitmapobjektet visas i mitten av sidan.  
Dra objektet till ett ställe där det är helt synligt, sedan upphäver du markeringen genom att klicka på något annat ställe.  
Objektet visas animerat.  
Redigera animerad GIF  
Om du vill redigera de enstaka bilderna i en animerad GIF-bild i efterhand, laddar du den animerade GIF-bilden till en sida i %PRODUCTNAME Impress och öppnar dialogrutan Animation (Bildskärmspresentation - Animation).  
Överta objekten med symbolen Överta objekt ett och ett.  
Radera nu alla bilder utom den önskade enstaka bilden och klicka på Skapa.  
Du kan sedan redigera denna enskilda bild på %PRODUCTNAME Impress-sidan.  
Därefter växlar du till den aktuella enstaka bilden i fönstret Animation, raderar den och övertar den markerade enskilda bilden från %PRODUCTNAME Impress-sidan.  
Spara animation som GIF-fil  
Markera objektet.  
Välj kommandot Arkiv - Exportera.  
Dialogrutan Exportera visas.  
Välj "GIF" (Graphics Interchange Format) som filtyp.  
Markera rutan Markering så att inte hela sidan exporteras, utan bara det markerade objektet.  
Välj en plats och ett namn för den animerade GIF-filen.  
Klicka på Spara.  
En animerad GIF-fil kan integreras i ett dokument på samma sätt som annan grafik (Infoga - Grafik).  
Du kan även använda Gallery för att ordna animerade GIF-bilder.  
Du behöver bara dra objektet från sidan till en temamapp i Gallery.  
Animera objekt till dia  
De effekter som används när du skiftar från en diabild till en annan kan du också använda vid visning av enskilda objekt eller objektgrupper.  
Vi vill visa en sida med en rubrik som "faller" på plats uppifrån.  
Därefter skall en rektangel glida in i bilden utmed en kurva som ritas fritt.  
1.  
Öppna ett nytt tomt presentationsdokument.  
2.  
Klicka på ikonen Text på verktygslisten, klicka sedan i dokumentet och skriv en text.  
Formatera texten om du vill.  
3.  
Välj kommandot Bildskärmspresentation - Effekt.  
Välj en effekt som på bilden ("Täck av uppifrån").  
4.  
Klicka på ikonen Tilldela.  
5.  
När du klickar i fönstret visas den aktuella effekten.  
Vid ett rent textobjekt (som alltså har skapats med verktyget Text, som i detta exempel) får symbolerna Effekter och Texteffekter samma resultat.  
Om du har en rektangel eller annat objekt, som du har dubbelklickat på och försett med en text, kan du däremot tilldela objektet och den tillhörande texten olika effekter.  
1.  
Rita nu en rektangel och ge den önskad färg.  
2.  
Rita en frihandslinje (utrullningslist Kurvor).  
3.  
Markera frihandslinjen och rektangeln (markeringsverktyg, håll ner skifttangenten).  
4.  
Välj Bildskärmspresentation - Effekt.  
5.  
I dialogrutan klickar du på Effekter.  
6.  
I listrutan väljer du "Övriga", sedan klickar du på Längs kurva.  
7.  
Klicka på Tilldela, och på Förhandsvisning om du vill.  
8.  
Om det finns flera objekt med effekter, kan du klicka på det objekt vars effekt du vill se i förhandsvisningen.  
9.  
Titta på presentationen genom att klicka på ikonen Bildskärmspresentation på verktygslisten.  
Om du har markerat rutan Manuell diabildsväxling i dialogrutan Bildskärmspresentation - Presentationsinställningar, måste du klicka med musen varje gång du vill växla diabild.  
I den här dialogrutan är varje effekt en "diabildsväxling".  
Animera diabildsväxling  
1.  
Skapa några sidor som innehåller objekt.  
Nya sidor skapar du t.ex. genom att klicka på det fria området till höger om sidflikarna vid arbetsområdets nedre kant.  
2.  
När du har ritat sidorna för en presentation byter du till diabildsvyn (Visa - Arbetsvy - Diabildsvy eller ikonen Diabildsvy i den högra kanten av fönstret).  
3.  
Du ser nu översikten över sidorna.  
Med ikonen Zoom kan du ändra skalan för översikten.  
4.  
Markera en dia och öppna dialogrutan Bildskärmspresentation - Diabildsväxling (eller Diabildsväxling på snabbmenyn till den markerade dian).  
Dialogrutan Diabildsväxling öppnas.  
I den här dialogrutan väljer du effekten som leder till att den markerade diabilden visas och som alltså syns innan diabilden är helt synlig.  
5.  
Du kan också välja effekter på diaobjektlisten där det finns olika listrutor, ikoner och rotationsfält där du kan ställa in effekter.  
Inställningarna som du gör här gäller direkt utan att du först måste klicka på Tilldela.  
6.  
Välj en effekt i den omfattande listan med effekter och klicka på Tilldela.  
Gör på samma sätt med de andra diabilderna som ska ha effekter.  
Om du klickar på den spelas en förhandsvisning av effekten upp på diabordet.  
Diabildsväxling  
Ordna dior på diabordet  
Växla till diabildsvyn.  
Ikonerna hittar du uppe till höger ovanför den högra rullningslisten.  
Här tilldelar du också effekterna för övergångarna.  
I diabildsvyn kan du dra diabilderna med musen och flytta dem till en annan plats så att diabildernas ordningsföljd ändras.  
Du kan kopiera en diabild med dra-och-släpp i diabildsvyn om du trycker på musknappen och Ctrl-tangenten och håller ner dem lite längre på diabilden.  
Muspekaren visar då ett plustecken.  
Det är också möjligt att använda dra-och-släpp från / till diabildsvyerna i andra %PRODUCTNAME Impress-dokument.  
Om du öppnar snabbmenyn till en markerad dia ser du också kommandot Visa diabild.  
Använd det här kommandot senare för att tillfälligt plocka ut den aktuella diabilden från din presentation, utan att radera den från dokumentet, för att sedan visa den igen.  
Namnet på en diabild som inte visas i presentationen markeras med grått i diabildsvyn.  
Arbetsvy  
Definiera bakgrundsfärg  
Bakgrunden på sidorna i ett tecknings - eller presentationsdokument kan du antingen rita och utforma i bakgrundsvyn eller så kan du tilldela sidorna en annan sidformatmall.  
Aktivera bakgrundsvyn med ikonen med samma namn i arbetsområdet nere till vänster.  
I bakgrundsvyn redigerar du bakgrunden för alla diabilder.  
Alla objekt, oavsett om det är företagslogotyper, linjer eller texter, som du matar in i den här vyn, visas i bakgrunden på alla sidor som använder den aktuella sidformatmallen (masterpage).  
På det här sättet kan du alltså reproducera sidhuvuden och sidfötter på presentationssidor.  
Objekten, som du infogar i bakgrundsvyn, är skyddade mot ändringar i normal sidvy.  
Det är också möjligt att ge bakgrunden en likformig struktur utan att bakgrundsvyn måste aktiveras:  
Välj Format - Sida och klicka på fliken Bakgrund i dialogrutan som visas.  
Välj ut en färg, färggradient, skraffering eller bitmap för bakgrunden.  
När du lämnar dialogrutan blir du tillfrågad om ändringen skall gälla för alla sidor eller bara för den aktuella sidan.  
Om du svarar med "Ja, ändringen skall gälla för alla sidor" ändras presentationsobjektmallen Bakgrund för den aktuella mastersidan.  
Alla diabilder som använder samma sidformatmall får den ändrade bakgrunden.  
Om du svarar med "Nej" ändras bara bakgrunden på den aktuella sidan.  
I %PRODUCTNAME Impress kan du också ändra presentationsobjektmallen i Stylist:  
Klicka på ikonen Presentationsobjektmallar i Stylist om den inte redan är intryckt.  
Du ser nu alla existerande mallar av den här typen i Stylist.  
Klicka på mallen Bakgrund.  
Öppna snabbmenyn till den här mallen och välj Ändra  
I dialogrutan som nu visas väljer du en passande färg till bakgrunden på alla sidor med den aktuella sidformatmallen.  
Klicka på OK.  
Den här ändringen av formatmallen gäller bara för det aktuella presentationsdokumentet.  
Ändra skala med tangent  
Om du vill förstora eller förminska vyn av ett grafikobjekt eller presentation eller återställa originalskalan kan du använda den numeriska delen av tangentbordet.  
Med minustangenten (-) förminskar du vyn, med plustangenten (+) förstorar du den.  
För varje gång du trycker på någon av tangenterna ändras skalan ett steg.  
Du återställer vyn till skala 1:1 med hjälp av tangenten bredvid minustangenten, på de flesta tangentbord har den ett multiplikationstecken (x)  
Kortkommandon för presentationer  
Exportera presentation som HTML  
Öppna presentationen som du vill exportera i HTML-format.  
Välj Arkiv - Exportera.  
Dialogrutan Exportera öppnas.  
Webbsida är redan valt som Filtyp.  
Ange ett Filnamn och klicka på Spara.  
AutoPilot för HTML-export öppnas.  
Den här AutoPiloten leder dig vidare med ett antal sidor.  
AutoPilot för HTML-export  
Arkiv - Exportera  
Importera HTML-sida till presentation  
Du kan importera en textsida, även i HTML-format, till en diabild från %PRODUCTNAME Impress.  
Växla till diabilden (till sidan) där textsidan eller HTML-sidan ska infogas.  
Välj Infoga - Fil.  
Dialogrutan Infoga fil öppnas.  
Du väljer "Text" eller "Webbsida "som Filtyp.  
Välj filen som ska infogas och klicka på Infoga.  
Om filen innehåller mer text än vad som får plats på en diabild fördelar du texten på flera diabilder:  
Klicka två gånger på den infogade texten så att du ser den gråa kanten som visar redigeringsläget.  
Markera all text som ligger nedanför den synliga diabilden och klipp ut den till urklippet - Kommando Ctrl +X.  
Infoga en ny tom diabild och klistra in innehållet från urklippet där - Kommando Ctrl +V.  
Upprepa de här stegen tills hela texten är fördelad på diabilderna.  
Individuell presentation  
Du kan visa dina diabilder från början till slut med t.ex. ikonen Bildskärmspresentation på verktygslisten eller med tangentkombinationen Kommando Ctrl +F2.  
I normala fall börjar en presentation alltid med den första diabilden.  
Om du alltid vill börja med den aktuella diabilden gör du så här:  
Välj Verktyg - Alternativ - Presentation - Allmänt.  
I området Starta presentation markerar du rutan Alltid med aktuell sida.  
Tänk på att den här inställningen har högre prioritet än den individuella presentationen som beskrivs nedan.  
Du har fler möjligheter att bara visa vissa diabilder eller att inte visa diabilder alls:  
Om du inte vill visa en dia väljer du diabildsvyn (t.ex. via menykommandot Visa - Arbetsvy - Diabildsvy), markerar diabilden och väljer Bildskärmspresentation - Visa diabild.  
Det signalerar att den inte visas i presentationen.  
Välj Bildskärmspresentation - Visa diabild när du vill visa diabilden igen.  
Du öppnar den på menyn Bildskärmspresentation.  
Klicka först på kommandoknappen Ny i dialogrutan Individuella bildskärmspresentationer.  
Dialogrutan Definiera individuell bildskärmspresentation öppnas.  
Här kan du ge presentationen ett namn.  
I den vänstra översikten över sidorna i presentationen markerar du en sida som du vill visa i den individuella presentationen och klickar på ikonen med pilen åt höger.  
Sidan infogas i det högra fältet.  
Alla sidor i det högra fältet visas i den individuella presentationen.  
Du kan arrangera om posterna i det högra fältet per dra-och-släpp med musen.  
Flytta objekt till annan nivå  
Om du vill flytta ett objekt från en nivå till en annan markerar du objektet och drar det till den andra nivåns registerflik.  
Låt musen vila ett ögonblick första gången Du har klickat och innan du flyttar muspekaren, så att objektet kan läggas till i urklippet.  
Infoga nivå  
Växla till nivåvyn, t.ex. med symbolen Nivåvy i symbolgruppen längst ned till vänster i arbetsområdet, eller via Visa - Nivå.  
I nedre kanten av arbetsområdet ser du registerflikarna för de fördefinierade nivåerna.  
Du kan visserligen använda de fördefinierade nivåerna, men inte döpa om eller radera dem.  
Klicka i det lediga området bredvid registerflikarna, eller välj kommandot Infoga nivå... i registerflikarnas snabbmeny.  
Dialogrutan Infoga nivå visas.  
Här ger du den nya nivån ett namn, och du kan också direkt bestämma om nivån ska vara synlig, utskrivbar eller spärrad.  
Klicka på OK.  
Den nya nivån är automatiskt den aktuella nivån, så att samtliga nu ritade objekt ligger på den nya nivån.  
Använda nivåer  
En del av dem kan du dölja, utesluta från utskrift eller spärra för fortsatt redigering.  
Nivåerna eller lagren är transparenta, vilket innebär att du alltid kan se alla nivåer samtidigt på alla sidor.  
Du kan göra varje enskild nivå osynlig och på detta sätt utesluta den från vyn.  
Du kan föreställa dig arbetet med nivåer som att alla dina objekt ligger ovanpå varandra på transparenta overheadblad.  
Det motsvarar visserligen inte helt nivåerna i %PRODUCTNAME, för nivåerna i %PRODUCTNAME definierar inte ordningsföljden mellan objekten när de ligger över varandra.  
Ordningsföljden mellan alla objekt i en stapel är snarare en egenskap som hör till varje enskilt objekt.  
Den är oberoende av den nivå där objekten finns.  
Varje sida i din teckning eller presentation kan innehålla flera nivåer, där det finns olika objekt.  
Men varje nivå existerar alltid samtidigt på alla sidor, och även bakgrunden kan innehålla flera nivåer.  
Tänk dig att du t.ex. gör planritningen till ett hus.  
På sidan 1 ritar du bottenvåningen, på sidan 2 vinden och på sidan 3 källaren.  
Väggarna med öppningar för dörrar och fönster ritar du enligt önskemål på grundnivån, d.v.s. på den nivå där du också ritar när du ännu inte vet något om nivåvyn (eller inte har aktiverat det).  
Denna nivå har namnet Layout.  
Alternativt kan du också definiera en ny nivå för väggarna med namnet "Väggar".  
Nu definierar du en nivå med namnet "Elektro" för elledningarna.  
Denna nivå gäller för samtliga sidor, men du kan placera olika objekt på nivån "Elektro" på varje sida.  
Naturligtvis kan nivån också vara helt tom på några sidor - eftersom alla nivåer är transparenta påverkar det inte synligheten för andra nivåer.  
På en annan nivå med namnet "Vatten" kan du rita in vattenledningarna.  
Nu kan du välja om du vill titta på och skriva ut alla nivåer för husets planritning, eller bara enstaka, eller valfria kombinationer.  
Men en nivå kan alltid bara vara synlig eller osynlig, utskrivbar eller inte utskrivbar för alla sidor gemensamt.  
Eftersom du först har ritat väggarna (oavsett på vilken nivå) och därefter elledningarna och vattenrören, ligger ledningarna och rören i objektstapeln över väggarna.  
Ordningsföljden i objektstapeln bestämmer du genom att markera ett eller flera objekt och sedan till exempel välja ikonerna på utrullningslisten Placering.  
Arbeta med nivåer  
Byta nivå  
Du byter till en annan nivå genom att växla till nivåvyn (Visa - Nivå) och sedan klicka på registerfliken för nivån.  
Dölja nivå  
Du kan snabbt göra en nivå synlig eller osynlig genom att hålla ner skifttangenten och klicka på registerfliken för nivån.  
Namnet på en osynlig nivå har blå färg.  
Spärra nivå  
Spärra en nivå om du vill se till att objekten på den nivån inte ändras mer.  
Om du ändå vill ändra dessa objekt måste du för säkerhets skull först upphäva spärren för nivån innan du kan ändra objekten eller lägga till nya objekt.  
Rita kurvor  
Verktygen för att rita kurvor och polygoner hittar du på utrullningslisten Kurvor.  
Dra listen till ett tomt tecknings - eller presentationsdokument.  
Klicka på ikonen Kurva.  
Markören blir till ett hårkors med en liten symbol som visar den nya funktionen.  
Nu kan du rita en kurva med nertryckt musknapp.  
Punkten där du först trycker på musknappen bestämmer startpunkten.  
Riktningen till den första punkten där du släpper musknappen, definierar riktningen som kurvan har från startpunkten.  
Nu flyttar du musen utan att trycka ner musknappen - kurvan följer musens rörelse - och klickar där den andra punkten i kurvan skall vara.  
Om du nu håller ner musknappen, kan du fortsätta (som när du hade tryckt första gången vid startpunkten) att bestämma kurvans riktning från den andra punkten till nästa, släppa musknappen och flytta musen vidare till punkt tre, klicka där igen och hålla ner musknappen och så vidare.  
Men om du släpper musknappen när du har klickat på kurvans andra punkt och sedan klickar på ett annat ställe på sidan, definierar du den andra punkten som hörnpunkt.  
I en hörnpunkt ändrar kurvan sin riktning abrupt med ett hörn.  
Om du även definierar punkt tre som hörnpunkt på det här sättet, får du en rät linje mellan punkt två och tre.  
Om du håller ner skifttangenten så är riktningarna begränsade till multipler av 45 grader.  
Om du håller ner Alternativ Alt -tangenten så sluts kurvan och du kan rita en annan kurva som kombineras med kurvan som precis slöts till ett gemensamt objekt.  
Om du vill sluta rita kurvor dubbelklickar du på den sista punkten som ska sättas.  
Du kan nu arbeta vidare med andra verktyg.  
De ritade kurvorna är Bézierkurvor.  
Punkterna på en Bézierkurva kallas för stödpunkter.  
Varje stödpunkt på Bézierkurvan kan vara "symmetrisk".  
Då har kurvan samma böjning på båda sidor om punkten.  
Då har kurvan olika böjningar på båda sidor av punkten.  
Om kurvan inte fortsätter i stödpunkten, utan har en hörna eller spets, rör det sig om en hörnpunkt.  
Du kan omvandla alla typerna till någon av de andra typerna och därmed utöva stort inflytande på kurvans form.  
Hur kan jag binda samman två punkter (t.ex. slutpunkter för linjer) exakt med linjer?  
För att exakt binda samman två punkter med linjer, använder du linjeikonen på verktygslisten.  
Dessutom måste alternativlisten vara aktiverad via Visa - Symbollister - Alternativlist.  
Aktivera ikonen Fäst mot objektpunkter på den här listen.  
Redigera kurva  
Du kan redigera stödpunkterna om de visas som små rektanglar.  
Om du vill redigera en kurva senare, när den inte längre är aktiverad, klickar du på ikonen Redigera punkter på Objektlisten och markerar kurvan.  
Om objektlisten inte är synlig klickar du kort på Urval på verktygslisten.  
Välj verktyget Redigera punkter längst till vänster på objektlisten eller på alternativlisten.  
Klicka en gång på punkten som du vill redigera.  
Den visas nu fylld och du ser båda stödlinjerna med kontrollpunkterna i ändarna.  
Vid hörnpunkter som definierar en rät vinkel ligger kontrollpunkterna direkt på stödpunkten.  
Du kan nu flytta stödpunkten och kontrollpunkterna fritt.  
Lägg märke till hur kurvan ändras motsvarande.  
Markören visar med sin respektive ändrade form vilken funktion du kan utföra.  
På objektlisten finns det några ikoner med vilka du bland annat kan ändra den markerade stödpunktens typ.  
En utförlig förklaring hittar du i %PRODUCTNAME -hjälpen.  
Om du vill omvandla typen av stödpunkt markerar du punkten.  
Hörnpunkt, Jämn övergång eller Symmetrisk övergång.  
Klicka på en ikon för den nya typen.  
Naturligtvis kan du också redigera kurvorna på "konventionellt vis", alltså ändra bredd, färg och vid fyllda kurvor även fyllningen.  
Alternativen för att ändra attributen hittar du på objektlisten när ikonen Redigera punkter inte är intryckt, på snabbmenyn och på menyerna Format och Ändra.  
Pröva även de andra ikonerna på utrullningslisten Kurvor.  
Om du avslutar en fylld kurva genom att dubbelklicka, sluts den automatiskt och sedan fylls alla "inre ytor".  
Objektlist  
Liveläge  
Tack vare det unika liveläget är det lätt att finputsa presentationer.  
En "riktig" presentation visas nog bara i helskärmsläge, därför är detta "standard ".  
Men för att redigera presentationen måste du egentligen växla till fönsterläge, så att du ser alla hjälpmedel, menyer och ikoner.  
I fönsterläget är proportionerna och helhetsintrycket helt annorlunda än i helskärmsläge.  
Liveläget löser det här problemet.  
Skapa eller öppna ett presentationsdokument.  
I det här exemplet räcker det även med en sida med ett enda objekt.  
Du gör inställningarna för typen av presentation med kommandot Bildskärmspresentation - Presentationsinställningar.  
De olika alternativen beskrivs utförligt i %PRODUCTNAME -hjälpen.  
Starta presentationen med standardinställningarna genom att klicka på ikonen Bildskärmspresentation på verktygslisten.  
När du ser den första diabilden (eller diabilden där du vill göra ändringar) öppnar du Navigator med F5.  
I Navigator klickar du på ikonen Liveläge.  
Nu kan du flytta, redigera och ändra alla objekt på sidan.  
Om du vill flytta objekt kan du bara ta tag i dem med musen och flytta dem.  
Andra egenskaper kan du ändra på snabbmenyn till det markerade objektet.  
Du ser ändringarna direkt i presentationen, i helskärmsläge.  
Stäng av liveläget i Navigator innan du avslutar presentationen.  
När liveläget är aktiverat kan du inte avsluta eller avbryta presentationen.  
Presentationsinställningar  
Anvisningar för %PRODUCTNAME Impress  
Göra och skriva ut presentation  
Animerade objekt och 3D-objekt  
Arbeta med nivåer  
Import och export  
Övrigt  
Byta sidformatmall  
Sidformatmallen bestämmer utseendet på objekten, inklusive bakgrunden, med sina underordnade formatmallar.  
Sidformatmallen kan också kallas för "masterpage".  
I %PRODUCTNAME Impress kan du tilldela varje sida en annan sidformatmall om du vill.  
Växla till sidan som skall få en annan masterpage.  
Välj Format - Formatmallar - Sidformatmall....  
Dialogrutan Sidformatmall visas.  
Dialogrutan Ladda sidformatmall visas.  
Välj en ny sidformatmall i dialogrutan, t.ex. i kategorin "Presentationsbakgrunder" och bekräfta med OK.  
Lägg märke till rutan Byt bakgrundssida.  
Om den inte är markerad gäller den nya sidformatmallen bara för den aktuella sidan.  
Du kan alltså tilldela en enskild sida en annan sidformatmall och därmed t.ex. en annan bakgrund.  
Den aktuella sidan får den nya bakgrunden som du har valt.  
Stylist  
Flytta objekt exakt på millimetern  
Om du vill flytta ett markerat objekt exakt horisontellt eller vertikalt använder du piltangenterna.  
Tryck på en av de fyra piltangenterna för att flytta objektet en millimeter.  
Utforma organisationsschema  
1.  
Du behöver för det första ett tomt teckningsdokument (Arkiv - Nytt - Teckning).  
2.  
Rita en tom eller en fylld rektangel med eller utan rundade hörn, som en namnskylt.  
Om du använder en fylld rektangel är det lättare att framhäva objekten med färg och det går att visa dem med skugga.  
3.  
För att alla namnskyltar skall bli lika stora duplicerar du den första namnskylten.  
Då är det ännu enklare att generera nästa namnskylt.  
Då kopieras inte bara nästa duplicerade namnskylt, utan även avståndet och riktningen till den föregående skylten kopieras.  
4.  
Ordna namnskyltarna bredvid respektive ovanför varandra så att de är centrerade.  
Välj sedan kommandot Justering - Centrerat på snabbmenyn eller på utrullningslisten Justering.  
5.  
När du har justerat namnskyltarna kan du skriva text på dem genom att dubbelklicka och sedan skriva texten.  
Du gör radbrytning med tangenterna Skift + Retur.  
6.  
Nu kan du förbinda två namnskyltar med varandra för att tydliggöra deras inbördes hierarkiska förhållande.  
Du väljer en typ av förbindelse mellan två namnskyltar på utrullingslisten Förbindelse.  
Om du nu pekar på en namnskylt (klicka inte ännu!) ser du hur skyltens kant blinkar.  
Det innebär att om du nu trycker på musknappen och drar musen till en annan namnskylt så har du fixerat förbindelsens första ankare vid hela objektet.  
Om du däremot pekar direkt på en av de fyra fördefinierade fästpunkterna mitt på objektets sidor, blinkar bara denna punkt.  
Drar du härifrån till ett annat objekt fästs förbindelsen vid denna punkt.  
Skillnaden mot den första metoden märker du när du flyttar ett objekt runt ett annat objekt.  
Om förbindelsen är fixerat vid hela objektet använder den alltid den fästpunkt som ligger närmast det andra objektet.  
När den andra metoden används stannar förbindelsen kvar vid den valda fästpunkten.  
Bestäm dig för en av metoderna och dra sedan musen från det ena objektet till det andra.  
Även vid målobjektet måste du destämma om du vill fixera förbindelsen vid en viss fästpunkt eller vid hela objektet.  
Vid cirklar, ellipser och 3D-objekt finns det fyra fördefinierade fästpunkter mitt på den begränsningsrektangelns sidor.  
Därför bör du själv definiera de önskade fästpunkterna vid sådana objekt.  
Du kan sedan välja om objektets fästpunkt skall ligga på kanten eller inne i objektet.  
1.  
När du ska placera en fästpunkt öppnar du alternativlisten (Visa - Symbollister - Alternativlist).  
Klicka på ikonen Redigera fästpunkter.  
Du ser nu fästpunktsobjektlisten (som du kan dra loss så att den blir ett eget fönster och senare förankra igen).  
2.  
Klicka på Infoga fästpunkt.  
Muspekaren visar sin nya funktion.  
3.  
Om inget objekt är markerat klickar du på ett objekt för att ange vilket objekt som ska få fästpunkten.  
Detta är nödvändigt eftersom fästpunkter även kan placeras utanför objektets yta (men de måste ligga innanför begränsningsrektangeln).  
4.  
Klicka på det ställe där du vill placera fästpunkten.  
Du ser där ett litet x.  
5.  
Du kan om du vill också låta förbindelser börja och sluta vid denna fästpunkt.  
Verktyget Infoga fästpunkt förblir aktiverat tills du väljer ett annat verktyg (t.ex. Urval).  
Du kan när som helst markera fästpunkter för att sedan flytta dem.  
Du kan också markera en förbindelse.  
Du kan också ändra typen, eller t.ex. ändra sträckningen i horisontell och vertikal riktning vid kurvförbindelser.  
Förbindelse  
Fästpunkter  
Kopiera sida från annan presentation  
Överföring av en sida från en presentation till en ny går till på följande sätt:  
Välj meny Infoga - Fil och välj ut den redan sparade presentationen.  
Om du trycker på kommandoknappen Infoga ser du en dialogruta som visar filen i trädstruktur.  
Om du klickar på ett plustecken, kan du välja ut och ladda den tillhörande sidan.  
Alternativt kan du välja sidan i diabildsvyn, kopiera den till urklippet och sedan klistra in den i det nya dokumentet.  
Infoga - Fil  
Ladda färgpaletter, färggradienter och skrafferingar  
Du sparar den aktuella färgpaletten och laddar en palett som fil med hjälp av symbolerna nere till höger under fliken Format - Yta - Färger.  
De leder till de vanliga dialogrutorna för val av filnamn och mappar.  
Som du ser om du tittar på de andra flikarna i dialogrutan Format - Yta kan du spara och ladda färggradienter, bitmapmönster och skrafferingar som fil.  
På detta sätt kan du skapa en passande omgivning för varje projekt.  
Du kan även ändra, spara och ladda linjestilar och linjeslut igen.  
Du redigerar dem i snabbmenyn för en linje.  
Du behöver alltså bara klicka på ikonen Spara i dialogrutan när du vill spara inställningarna med ett annat namn.  
%PRODUCTNAME levereras med många alternativa färgpaletter, färggradienter, skrafferingar, linjestilar och linjeslut.  
De här objekten finns i filerna i mappen {installpath} / user / config.  
I förinställningen är alltid filen "Standard" öppen.  
I filerna med namnen "Standard" är namnen på de medföljande objekten på engelska, men de översätts internt beroende på din språkversion av %PRODUCTNAME.  
Därigenom garanteras en språkövergripande användning av dessa objekt.  
Typ  
Ändelse  
Exempel  
Färgpaletter  
*.soc  
CMYK, palett, webb, HTML, standard  
Färggradienter  
*.sog  
classic, modern, standard  
Skrafferingar  
*.soh  
Skraffering, standard  
Linjestilar  
*.sod  
Stilar, standard  
Linjeslut  
*.soe  
Slut, standard  
Lägg särskilt märke till färgpaletten Cmyk.soc som hjälper dig att optimalt återge färgglad grafik i CMYK-kulörsystem på papper.  
Färgpaletten Web.soc innehåller en särskild World Wide Web-färgpalett med 16 standardfärger och 216 RGB-färger uppbyggda efter ett visst schema.  
Färgpaletten HTML.soc har ett liknande användningsområde.  
Du kan titta på några färgpaletter i %PRODUCTNAME Draw-exempeldokumentet "Färgprofil".  
I det här dokumentet finns även %PRODUCTNAME -standardfärgerna.  
Format - Yta  
Skriva ut presentationer  
Välja förinställningar för alla utskriftsjobb  
Klicka på Presentation - Skriv ut.  
Inställningarna som du gör här gäller för alla utskriftsjobb.  
Välja utskriftsalternativ för den aktuella utskriften  
Välj kommandot Arkiv - Skriv ut.  
Dialogrutan Skriv ut öppnas.  
Klicka på Fler.  
Dialogrutan Skrivaralternativ.  
Inställningarna i den här dialogrutan gäller bara för det aktuella utskriftsjobbet.  
Skriva ut anteckningar, flygblad, disposition  
Välj utskriftsalternativ enligt beskrivningen ovan, antingen för alla utskriftsjobb eller för den aktuella utskriften.  
Skriva ut utvalda diabilder  
Växla till diabildsvyn, t.ex. med ikonen Diabildsvy på den högra rullningslisten.  
Håll ner skifttangenten och klicka på alla diabilder som du vill skriva ut.  
Diabilderna får en markering i kanten.  
Välj kommandot Arkiv - Skriv ut.  
Dialogrutan Skriv ut öppnas.  
De markerade sidorna = diabilderna är angivna som Utskriftsområde.  
Klicka på OK.  
Anpassa utskrift till papperssida  
Kan ett dokument som är skapat i format A0 skrivas ut i A4-storlek?  
Om du vill förminska en sida i %PRODUCTNAME Draw / %PRODUCTNAME Impress till t.ex. A4-format med rätt proportioner, måste den här anpassningen väljas vid inställningen av sidan.  
1.  
Ladda ditt dokument med A0-sidan.  
2.Välj Sida - Ställ in sida på snabbmenyn.  
3.  
I dialogrutan markerar du rutan Anpassa objekt till pappersformat i området Layoutinställningar.  
4.  
Ändra sidstorleken till A4 och anpassa ev. sidans marginaler.  
5.  
Klicka på OK.  
De relativa positionerna är desamma.  
Du kan också välja att skriva ut direkt.  
Då visas en dialogruta som frågar dig om sidan skall anpassas till utskriftsområdet, skrivas ut på flera sidor eller kortas av.  
Markera täckt objekt  
Om du vill markera ett objekt som är helt täckt av ett annat objekt håller du ner Alternativ Alt -tangenten och klickar på objektets plats.  
Om du dessutom håller ner skifttangenten går du igenom objekten i andra riktningen varje gång du klickar.  
Du markerar ett objekt med tabbtangenten.  
Nästa objekt markeras när du trycker på tabbtangenten igen.  
Med Skift-Tabb byter du riktning bland objekten.  
Infoga tabell på diabild  
Infoga en ny tabell  
Växla till diabilden där du vill skriva om tabellen.  
Välj en sidlayout med tabell:  
Välj Format - Ändra sidlayout.  
Dubbelklicka på autolayouten med namnet Rubrik, tabell.  
Dubbelklicka på platshållaren för tabellen.  
Du kan mata in data, formatera celler, klistra in innehåll.  
Klicka utanför tabellen för att avsluta inmatningen.  
Klicka en gång på tabellen om du vill flytta, radera eller skala den.  
Dubbelklicka på tabellen för att redigera den.  
Infoga ett %PRODUCTNAME Calc-dokument  
Växla till diabilden där du vill infoga tabellen i form av ett dokument.  
Välj kommandot Infoga - Objekt - OLE-objekt.  
Dialogrutan Infoga OLE-objekt öppnas.  
Välj alternativet Skapa från fil.  
Klicka på Genomsök och välj ut det önskade dokumentet.  
Format - Ändra sidlayout  
Infoga - Objekt - OLE-objekt  
Omvandla texttecken till kurvor  
Skriv texten eller bokstaven resp. specialtecknet i ett %PRODUCTNAME Draw-dokument.  
Välj en lämplig teckenstorlek och ett lämpligt teckensnitt.  
Om du vill skriva text klickar du på ikonen Text på utrullningslisten Text från verktygslisten.  
Låt textobjektet vara markerat och välj Ändra - Omvandla - Till kurva.  
Texten omvandlas till en Bézierkurva.  
Om texten består av mer än ett tecken har du nu en grupp av objekt.  
För att kunna redigera ett enskilt tecken går du in i grupperingen.  
Välj t.ex. Gå in i gruppering på snabbmenyn till gruppen eller tryck på F3.  
Klicka därefter på tecknet som du vill redigera.  
Klicka på ikonen Redigera punkter (uppe till vänster på bilden).  
Klicka på objektet.  
På objektlisten finns ikonerna för redigering, infogning och radering av punkterna.  
Använd utrullningslisten Zoom för att förstora vyn.  
Om skrivtecknens svarta fyllning stör vid redigeringen ändrar du den tillfälligt till t.ex. 10% grått med kommandot Format - Yta.  
Format - Yta  
Vektorisering av en bitmap  
Du kan också omvandla pixelbilder, såkallade bitmaps, till vektorteckningar med %PRODUCTNAME Impress eller %PRODUCTNAME Draw.  
Vektorgrafikobjekt har bland annat den fördelen att de ser bra ut vid utskrift oavsett vilken skala de har.  
Vid utskrift av skalade bitmaps förekommer det ofta fula trappeffekter, grova klossraster eller att fina linjer saknas.  
1.  
Välj den bitmap som du vill vektorisera, t.ex. genom att klicka en gång på objektet.  
2.  
Välj Omvandla - Till polygon.  
I %PRODUCTNAME Draw hittar du kommandot under meny Ändra, i %PRODUCTNAME Impress på snabbmenyn till det markerade objektet.  
Du ser dialogrutan Omvandla till polygon.  
Här kan du ställa in några parametrar för omvandlingen och se en förhandsvisning av resultatet.  
3.  
Om du klickar på OK ersätts den markerade bitmappen med ett vektorgrafikobjekt som metafil.  
Välkommen till %PRODUCTNAME Impress-hjälpen  
Hjälp till %PRODUCTNAME Impress  
Hjälp till hjälpen  
Menyer  
Här hittar du beskrivningen av alla menyer med undermenyer och dialoger.  
Arkiv  
I den här menyn finns kommandon för hantering av dokument som helhet.  
Du kan t.ex. skapa ett nytt dokument, öppna, stänga, och skriva ut dokument, ange dokumentegenskaper med mera.  
När du vill avsluta %PRODUCTNAME Impress klickar du på menykommandot Avsluta.  
Öppna...  
Spara som...  
Exportera...  
Versioner...  
Egenskaper...  
Skriv ut...  
Skrivarinställning...  
Redigera  
Här finns bl.a. kommandona som du använder när du vill ångra den senaste åtgärden, kopiera och klistra in via urklippet och öppna dialogrutan Sök och ersätt.  
Klistra in innehåll...  
Sök och ersätt...  
Duplicera...  
Fältkommando...  
Radera sida...  
Länkar...  
Image map  
Hyperlänk  
Visa  
Den här menyn innehåller kommandon som används till styra hur dokumentinnehållet ser ut på bildskärmen.  
Skala...  
Infoga  
På den här menyn är alla kommandon sammanfattade som används till att infoga nya element i dokumentet, som t.ex. skannade objekt, grafik, objekt, symboler och andra filer.  
Sida...  
Specialtecken...  
Hyperlänk  
Tabell  
Ritobjekt som har infogats på ritbordet centreras inte på sidan.  
Diagram...  
Ram...  
Fil...  
Format  
Här hittar du kommandona som används till att ställa in objekt - och sidformateringen.  
Vid markerade objekt ändras menyn och deras speciella formatkommandon visas.  
I den här menyn hittar du dessutom funktionerna för hantering av mallar, t.ex. mallkatalogen och Stylist.  
Linje...  
Yta...  
Text...  
Position och storlek...  
Kontrollfält...  
Formulär...  
Dimensionering  
Förbindelse...  
Tecken...  
Numrering / punktuppställning...  
Stycke...  
Sida...  
Ändra sidlayout...  
Verktyg  
Menyn Verktyg innehåller kommandon beträffande lingvistik och diverse programalternativ.  
Här startar du rättstavningskontrollen eller synonymordlistan som kan föreslå alternativ till ord.  
Dessutom kan du anpassa utseendet på symbollister och menyer, konfigurera tangentbordet och göra allmänna standardinställningar för programmet.  
Synonymordlista...  
AutoKorrigering...  
Makro...  
Anpassa...  
Fönster  
I fönstermenyn kan du öppna fönster.  
Där finns också en lista över öppna dokument.  
Ändra  
Den här menyn innehåller kommandon för att redigera objekt, som t.ex. Spegelvänd, Omvandla till kurvor, Placering och Justering.  
Fördelning...  
Namnge objekt...  
Gruppering  
Upphäv gruppering  
Gå in i gruppering  
Lämna gruppering  
Bildskärmspresentation  
I den här menyn har du många olika möjligheter att utforma presentationens förlopp på ett optimalt sätt.  
Presentationsinställningar...  
Individuell bildskärmspresentation...  
Interaktion...  
Symbollister  
Här hittar du en beskrivning av elementen på symbollisterna i ett aktivt presentationsdokument.  
Objektlist teckningsvy, anteckningsvy, flygbladsvy  
På den här objektlisten hittar du funktionerna som du behöver i det aktuella redigeringsläget.  
Linjestil  
Linjebredd  
Linjefärg  
Ytstil - / fyllning  
Skugga  
Objektlist vid textinmatning  
Objektlisten visas när textmarkören står i texten.  
Det finns två objektlister för textredigering som skiljer sig något åt.  
I den högra kanten av objektlisten finns det en liten svart trekant för att växla mellan den och alla andra aktiva objektlister.  
Med följande ikoner formaterar du texten direkt, utan formatmallar.  
Med kommandot Format - Standard kan du ta bort alla direkta formateringar i den markerade texten.  
Teckenfärg  
Tecken  
Stycke  
Punktuppställningstecken  
Objektlist i diabildsvyn  
På objektlisten i diabildsvyn i %PRODUCTNAME Impress kan du bl.a. välja toningseffekter mellan diabilderna.  
På verktygslisten i diabildsvyn finns dessutom ett zoomnings - och ett urvalsverktyg med vars hjälp du kan titta på sidorna i presentationen och sortera dem genom att dra och släppa dem.  
Statuslist  
Där finns även några kommandoknappar med specialfunktioner.  
Linjaler  
Linjalerna i den vänstra och övre kanten av fönstret i ett %PRODUCTNAME Impress-dokument visar hela tiden sidans mått samt det aktuella objektets placering och storlek.  
Du kan visa eller dölja linjalerna med kommandot Visa - Linjaler.  
Den öppnar du genom att placera muspekaren på en av linjalerna, hålla ner Ctrl-tangenten och klicka med högra musknappen.  
Du kan läsa av måtten för ett markerat objekt direkt på markeringarna på linjalerna.  
Om du drar i en sådan markering med musen ändras objektets storlek.  
Du kan även ändra sidmarginalerna genom att dra i kanterna på det vita området på linjalerna.  
Om du vill flytta nollpunkten för koordinaterna som visas kan du dra skärningspunkten för de båda linjalerna uppe till vänster till önskat läge (som dock måste ligga innanför sidmarginalerna).  
Om du dubbelklickar här flyttas nollpunkten till sidans övre vänstra hörn.  
Om du drar med musen från linjalområdet till sidan kan du infoga ett valfritt antal stödlinjer, som objekten fäster mot vid flyttning eller storleksförändring.  
När du redigerar ett textobjekt visas tabbarna på linjalen och kan ändras där.  
Verktygslisten i tecknings-, antecknings - och flygbladsvyn  
Enligt standardinställningen visas den här verktygslisten till vänster om dokumentet.  
På den här förankringsbara listen är de viktigaste redigeringsfunktionerna tillgängliga.  
Flera av ikonerna är utrullningslister, som i sin tur innehåller fler ikoner.  
Ikonerna med utrullningslister är markerade med små trekanter.  
Markera objekt  
Du kan markera objekt genom att klicka på dem med urvalsverktyget.  
Om du håller ner skifttangenten när du klickar kan du markera flera objekt samtidigt.  
Om flera objekt ligger staplade på varandra kan du markera dolda objekt genom att hålla ner Alternativ Alt -tangenten när du klickar.  
Om du håller ner Skift + Alternativ Alt -tangenten markeras föregående objekt i stapeln nästa gång du klickar.  
De flesta redigeringsverktygen påverkar objekt som är markerade.  
Ett markerat objekt har åtta små handtag.  
Om du dubbelklickar på ett markerat objekt kan du mata in en text som är kopplad till objektet.  
Upphäv markeringen genom att klicka utanför det markerade objektet.  
Rotera  
Med det här verktyget kan du rotera ett objekt.  
Det motsvarar kommandot Rotera, som även finns på verktygslisten i %PRODUCTNAME Draw under Effekter.  
Interaktion  
Verktygslisten i dispositionsvyn  
Enligt standardinställningen visas den här verktygslisten till vänster om dokumentet när du har aktiverat dispositionsvyn i menyn Visa - Arbetsvy.  
På den här förankringsbara listen finns de viktigaste redigeringsfunktionerna.  
En del av ikonerna är utrullningslister som i sin tur innehåller andra ikoner.  
Ikonerna med utrullningslister är markerade med små trekanter.  
Bildskärmspresentation  
Verktygslisten i diabildsvyn  
Enligt standardinställningen finns den här verktygslisten till vänster om dokumentet när du har aktiverat diabildsvyn i menyn Visa - Arbetsvy.  
På denna förankringsbara list finns de viktigaste redigeringsalternativen.  
Vissa av ikonerna är utrullningslister som i sin tur innehåller andra ikoner.  
Ikonerna med utrullningslister är markerade med en liten trekant.  
Bildskärmspresentation  
Alternativlist  
På den här förankringsbara listen har du tillgång till viktiga alternativ utan att behöva öppna enskilda dialogrutor.  
Visa raster  
Hjälplinjer vid förflyttning  
Fäst mot raster  
Fäst mot stödlinjer  
Fäst mot sidmarginaler  
Fäst mot objektram  
Fäst mot objektpunkter  
Tillåt snabbredigering  
Bara textområde kan markeras  
Antyd extern grafik  
Konturläge  
Antyd text  
Visa bara fina linjer  
Grafikobjektlist  
Om ett grafikobjekt är markerat i ett dokument visas grafikobjektlisten.  
Funktioner i %PRODUCTNAME Impress  
Här får du en kort överblick över några viktiga funktioner i %PRODUCTNAME Impress.  
För kontorsanvändare ger %PRODUCTNAME Impress bra hjälp.  
Utforma vektorgrafik  
I %PRODUCTNAME Impress har du tillgång till nästan alla verktyg som också finns i %PRODUCTNAME Draw när du ska utforma vektorgrafik.  
Diabildsvisning  
%PRODUCTNAME Impress kan hantera nästan hur många sidor som helst i ett enskilt dokument.  
Varje sida motsvarar en dia - eller OH-bild i en presentation.  
Mallkonceptet i %PRODUCTNAME gör det enkelt för dig att ge alla dina diabilder ett enhetligt utseende.  
Bildspelen i %PRODUCTNAME Impress kan lättas upp med hjälp av ett stort antal effekter.  
Du kan lägga in en ljudeffekt eller tilldela objekten på varje sida en animation och en effekt som du aktiverar genom att klicka på objektet med musen.  
Utveckla presentationer  
Det finns fler hjälpmedel i %PRODUCTNAME Impress när du skapar presentationer.  
Du kan växla till dispositionsvyn för att ordna och strukturera dina idéer.  
I diabildsvyn ser du en översikt av diabilderna och kan gruppera om, kopiera, klippa ut och infoga dem även utanför det synliga området genom att dra och släppa.  
I flygbladsvyn kan du skriva ut åhörarkopior.  
Om du provkör presentationen kan du använda automatisk tidtagning och lägga in den tid som t.ex. behövs för det du ska säga för varje enskild dia.  
Publicera presentationer  
Exportera din presentation med hjälp av en speciell AutoPilot så att du kan publicera den på Internet.  
Alla konverteringar som är nödvändiga utförs automatiskt.  
Den exporterade presentationen kan visas med alla moderna webbläsare.  
Framföra livepresentationer  
Under presentationens gång kan du rita på diabilderna med musen för att betona viktiga punkter, precis som med en markeringspenna.  
I liveläget kan du ändra och radera objekt på diabilderna och lägga till nya objekt medan presentationen pågår.  
Så hittar du den här funktionen...  
Menyn Redigera - Nästa platshållare  
Tangenten F2  
Menyn Redigera - Föregående platshållare  
Tangentkombinationen Skift+F2  
Menyn Redigera - Nästa fel  
Tangenten F3  
Menyn Redigera - Föregående fel  
Tangentkombinationen Skift+F3  
Ikon på verktygslisten:  
Zoom 100%  
Menyn Visa - Förstora  
Ikon på verktygslisten:  
Större  
Menyn Visa - Förminska  
Ikon på verktygslisten:  
Mindre  
Menyn Visa - Visa allt  
Ikon på verktygslisten:  
Hela formeln  
Menyn Visa - Uppdatera  
Tangenten F9  
Ikon på verktygslisten:  
Uppdatera  
Menyn Visa - Uppdatera visning automatiskt  
Menyn Visa - Urval  
Snabbmenyn i kommandofönstret - Monära / Binära operatorer  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Unära / Binära operatorer  
Snabbmenyn i kommandofönstret - Relationer  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Relationer  
Snabbmenyn i kommandofönstret - Operatorer  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Operatorer  
Snabbmenyn i kommandofönstret - Funktioner  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Funktioner  
Snabbmenyn i kommandofönstret - Parenteser  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Parenteser  
Snabbmenyn i kommandofönstret - Attribut  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Attribut  
Snabbmenyn i kommandofönstret - Formateringar  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Formateringar  
Snabbmenyn i kommandofönstret - MÃ¤ngdoperationer  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Mängdoperationer  
Menyn Format - Teckensnitt...  
Menyn Format - Teckensnitt - Ã„ndra -...  
Menyn Format - Teckenstorlekar...  
Menyn Format - AvstÃ¥nd...  
Menyn Format - Justering...  
Menyn Format - TextlÃ¤ge  
Menyn Verktyg - Katalog  
Ikon på verktygslisten:  
Symboler  
Menyn Verktyg - Katalog - Redigera  
Menyn Verktyg - Importera formel...  
Menyn Verktyg - Anpassa  
Snabbmenyn i kommandofönstret - Övrigt  
Menyn Visa - Urval - ikon i urvalsfönstret:  
Övrigt  
Formelmarkör  
Nästa platshållare  
Sätter markören på nästa platshållare.  
Platshållare visas i form av <?> i fönstret Kommandon.  
Föregående platshållare  
Sätter markören på den föregående platshållaren.  
Platshållare visas i form av <?> i fönstret Kommandon.  
Nästa fel  
Placerar markören på nästa fel  
Föregående fel  
Placerar markören på det föregående felet.  
Förstora  
Skalan förstoras med 25%.  
Skalan visas på statuslisten.  
Du kan även ändra skalan på snabbmenyn där.  
Även snabbmenyn i arbetsområdet innehåller en urvalslista.  
Förminska  
Skalan förminskas med 25%.  
Skalan visas på statuslisten.  
Du kan även ändra skalan på snabbmenyn där.  
Även snabbmenyn i arbetsområdet innehåller en urvalslista.  
Visa allt  
Här ställer du in visningen så att du ser hela formeln i maximal storlek.  
Formeln förminskas eller förstoras i arbetsområdet så att alla formelelement syns.  
Visa allt motsvarar ikonen Hela formeln på verktygslisten.  
På statuslisten visas den för tillfället aktuella skalan.  
Om du öppnar snabbmenyn där, så visas en urvalslista med tillgängliga skalor för visningen.  
Även med snabbmenyn för arbetsområdet kan du öppna en urvalslista.  
Uppdatera  
Med det här kommandot ritar du om formeln i dokumentfönstret.  
Ändringar som du gör i fönstret Kommandon uppdateras automatiskt om Uppdatera visning automatiskt är aktiverat.  
Uppdatera visning automatiskt  
Aktivera det här kommandot om du vill att en ändrad formel ska uppdateras automatiskt.  
Om du inte väljer det här alternativet, ritas formeln först om med kommandot Visa - Uppdatera (F9).  
Urval  
Här finns ikoner som du använder när du ska infoga operatorer, funktioner, symboler och ändra layout.  
Några exempel visar vilka funktioner som finns.  
Det finns fler exempel för formeldokument i mappen Exempel - Formler.  
Urvalsfönstret är indelat i två områden.  
Om du klickar på en ikon i det övre området visas de tillhörande ikonerna i det undre området.  
I fönstret Kommandon visas det indelade urvalet som undermenyer.  
Referens  
Unära / binära operatorer  
Välj bland de olika unära och binära operatorerna till din %PRODUCTNAME Math -formel.  
Unära operatorer verkar på "en" platshållare, medan binära sätter "två "platshållare i relation till varandra.  
De olika operatorerna visas i det undre området i urvalsfönstret.  
Du kan även visa en lista över samma funktioner och några fler genom att öppna snabbmeny n i fönstret Kommandon.  
Alla operatorer som inte finns med i urvalsfönstret måste du ange direkt i kommandofönstret.  
Du kan göra alla infogningar direkt, även dem för vilka det finns ikoner.  
Operatorer som listas tillsammans med en ikon kan du infoga via urvalsfönstret (menyn Visa - Urval) och snabbmenyn (kommandofönstret).  
De olika unära och binära operatorerna är:  
Tecken +  
Med den här ikonen infogar du ett plustecken med platshållare.  
Tecken -  
Med den här ikonen infogar du ett minustecken med platshållare.  
Skriv sedan - <?> i kommandofönstret.  
Tecken plus / minustecken  
Med den här ikonen infogar du ett plus / minustecken med platshållare.  
Du kan skriva den här operatorn direkt i kommandofönstret genom att först skriva plustecknet, sedan minustecknet och till slut platshållaren.  
Minus / plustecken  
Med den här ikonen infogar du ett minus / plustecken med platshållare.  
Du kan skriva den här operatorn direkt i kommandofönstret genom att först skriva minustecknet, sedan plustecknet och till slut platshållaren.  
Addition  
Med den här ikonen infogar du en addition med två platshållare.  
I kommandofönstret kan du i stället ange <?> + <?>.  
Multiplikation (punkt)  
Multiplikation; tecken som punkt Med den här ikonen infogar du en multiplikation med en liten multiplikationspunkt och två platshållare.  
Du kan också skriva <?>cdot<?> i kommandofönstret.  
Multiplikation (x)  
Med den här ikonen infogar du en multiplikation med två platshållare.  
Som multiplikationstecken används ett kryss.  
Du kan också skriva <?>times<?> i kommandofönstret.  
Multiplikation (*)  
Med den här ikonen infogar du en multiplikation med två platshållare.  
Som multiplikationstecken används här en asterisk.  
Du kan också skriva <?> * <?> i kommandofönstret.  
Tecken + -  
Med den här ikonen infogar du en subtraktion med två platshållare.  
Du kan också skriva <?> - <?> i kommandofönstret.  
Division (bråk)  
Med den här ikonen infogar du ett bråk med två platshållare.  
Du kan också skriva <?> over <?> direkt i kommandofönstret.  
Division (kolon / snedstreck)  
Med den här ikonen infogar du en division med två platshållare.  
Du kan också skriva <?> div <?> i kommandofönstret.  
Division (snedstreck)  
Med den här ikonen infogar du en division med två platshållare.  
Men som divisionstecken används ett snedstreck /.  
Du kan också skriva <?> / <?> i kommandofönstret.  
Logiskt INTE  
Med den här ikonen infogar du tecknet för ett logiskt INTE med platshållare.  
Du kan också skriva neg <?> direkt i kommandofönstret.  
Logiskt OCH  
Med den här ikonen infogar du en logisk OCH-operator.  
Du kan också skriva <?> and <?> i kommandofönstret..  
Logiskt ELLER  
Med den här ikonen infogar du en logisk ELLER-operator.  
Du kan också skriva <?> or <?> i kommandofönstret.  
Länkning  
Med den här ikonen infogar du en länkning av symboler.  
Du kan också skriva circ i kommandofönstret.  
Det är bl.a. särskilt användbart om du vill bygga in speciella tecken i en formel.  
Den här typen av operator använder du enligt följande mönster: uoper %theta x.  
Som exempel skapas här den lilla grekiska bokstaven theta, som ingår i %PRODUCTNAME Math -teckenuppsättningen.  
Du kan även använda operatorn om du vill infoga tecken som inte kommer från %PRODUCTNAME.  
Men då måste du först göra det önskade tecknet tillgängligt via menyn Verktyg - Symboler - Katalog... - Redigera.  
Med boper kan du infoga användardefinierade binära operatorer.  
Det är bl.a. särskilt användbart om du vill bygga in speciella tecken i en formel.  
Den här typen av operator använder du enligt följande mönster: x boper %theta y.  
I exemplet skapas den lilla grekiska bokstaven theta.  
Den här operatorn är särskilt intressant eftersom du kan använda den när du vill infoga tecken som inte kommer från %PRODUCTNAME.  
Även för den här operatorn måste du först göra motsvarande inställningar i menyn Verktyg - Symboler.  
Med kommandot <?>oplus<?> infogar du ett additionstecken som omges av en cirkel i dokumentet.  
Med <?>ominus<?> infogar du ett subtraktionstecken som omges av en cirkel.  
Genom att skriva <?>odot<?> i kommandofönstret infogar du en multiplikationspunkt i en cirkel.  
Med <?>odivide<?> infogar du ett snett divisionsstreck som omges av en cirkel i formeldokumentet.  
Med kommandot a wideslash b skapar du två tecken med ett mellanliggande diagonalt streck som börjar nerifrån vänster och sträcker sig uppåt åt höger.  
Tecknens höjd justeras så att tecknet till vänster om strecket höjs och tecknet till höger sänks.  
Det här kommandot når du även via kommandofönstrets snabbmeny, men inte via urvalsfönstret.  
Med kommandot a widebslash b infogar du två tecken med ett mellanliggande diagonalt streck som börjar nerifrån höger och sträcker sig upp till vänster.  
Tecknens höjd justeras så att tecknet till vänster om strecket sänks och tecknet till höger höjs.  
Det här kommandot når du även via kommandofönstrets snabbmeny, men inte via urvalsfönstret.  
Kommandona sub och sup kan du använda för att lägga till index och potenser till tecknen i formeln, t.ex. a sub 2.  
Vill du använda kolon (:) som divisionstecken?  
Då öppnar du dialogrutan Symboler via menyn Verktyg - Symboler - Katalog....  
Du kan även öppna den här dialogrutan via ikonen på verktygslisten.  
Klicka sedan på kommandoknappen Redigera....  
Dialogrutan Redigera symboler öppnas.  
Ange ett så beskrivande namn som möjligt i kombinationsfältet Symbol, t.ex. delad, och klicka på det önskade tecknet i symbolsetets visningsfält.  
Klicka först på kommandoknappen Lägg till och sedan på OK.  
Stäng dialogrutan Symboler med Stäng.  
Nu kan du använda den nya symbolen enligt mönstret a %delad b = c.  
När du skriver in något manuellt i kommandofönstret bör du tänka på att blankstegen är absolut nödvändiga för att du ska åstadkomma korrekt uppbyggnad för många operatorer.  
Detta gäller i synnerhet om du förser operatorerna med värden i stället för med platshållare, t.ex. om du bygger upp divisionen 4 div 3 eller a div b.  
Relationer  
Välj den relation som du vill använda i din %PRODUCTNAME Math -formel.  
Alla relationer som är tillgängliga i urvalsfönstret hittar du i det undre området i fönstret.  
En motsvarande lista visas även om du öppnar snabbmeny n i fönstret Kommandon.  
Relationer som du inte kan nå via urvalsfönstret måste du skriva in direkt i kommandofönstret.  
Alla infogningar för vilka det finns ikoner kan du givetvis även göra manuellt.  
Det är bara relationer som listas tillsammans med en ikon som du kan infoga via urvalsfönstret (menyn Visa - Urval) och snabbmenyn (kommandofönstret).  
De olika relationerna är:  
är lika med  
Med den här ikonen infogar du ett likhetstecken med två platshållare.  
Du kan också skriva <?> = <?> i kommandofönstret.  
är inte lika med  
Med den här ikonen eller med kommandot neq infogar du en olikhet med två platshållare.  
I stället för neq kan du använda tecknen <>.  
Du gör inmatningen enligt mönstret <?>neq<?>.  
är kongruent med  
Med den här ikonen infogar du ett tecken för relationen kongruent med två platshållare.  
Du kan också skriva <?>equiv<?> i kommandofönstret.  
är ortogonal med  
Med den här ikonen infogar du ett tecken för en rätvinklig (ortogonal) relation med två platshållare.  
Du kan också skriva <?>ortho<?> direkt i kommandofönstret.  
delar  
Med den här ikonen infogar du tecknet för "delar".  
Du kan också skriva <?> divides <?> i kommandofönstret.  
delar ej  
Med den här ikonen infogar du tecknet för "delar ej".  
Du kan också skriva <?> ndivides <?> i kommandofönstret.  
är mindre än  
Med den här ikonen infogar du relationen "mindre än".  
I ställte för att använda ikonen kan du skriva <?> lt <?> eller < i kommandofönstret.  
är större än  
Med den här ikonen infogar du relationen "större än".  
I stället för att använda ikonen kan du skriva <?> gt <?> eller > i kommandofönstret.  
är ungefär lika med  
Med den här ikonen infogar du ett tecken för relationen ungefär med två platshållare i dokumentet.  
Du kan även skriva <?>approx<?> direkt i kommandofönstret.  
är parallell med  
Med den här ikonen infogar du en parallell relation med två platshållare.  
Du kan också skriva <?>parallel<?> direkt i kommandofönstret.  
är mindre än eller lika med (sned)  
Med den här ikonen infogar du relationen "är mindre än eller lika med" med två platshållare.  
Du kan även skriva <?>leslant<?> direkt i kommandofönstret.  
är större än eller lika med (sned)  
Med den här ikonen infogar du relationen "är större än eller lika med" med två platshållare.  
Du kan även skriva <?>geslant<?> direkt i kommandofönstret.  
är liknande eller lika med  
Med den här ikonen infogar du en "är liknande eller lika med "-relation med två platshållare.  
Du kan också skriva <?>simeq<?> direkt i kommandofönstret.  
är proportionell mot  
Med den här ikonen infogar du relationen "är proportionell mot" med två platshållare.  
Du kan också skriva <?>prop<?> direkt i kommandofönstret.  
är mindre än eller lika med  
Med den här ikonen infogar du relationen "mindre än eller lika med" med två platshållare.  
Du kan också skriva <?> le <?> eller <= direkt i kommandofönstret.  
är större än eller lika med  
Med den här ikonen infogar du relationen "större än eller lika med" med två platshållare.  
I stället för att använda ikonen kan du skriva <?>ge<?> eller >=.  
liknar  
Med den här ikonen infogar du relationen "liknar" med två platshållare.  
Du kan också skriva <?>sim<?> i kommandofönstret.  
strävar mot  
Med den här ikonen infogar du relationen "strävar mot" med två platshållare.  
Du kan också skriva <?>toward<?> i kommandofönstret.  
dubbelpil till vänster  
Med den här ikonen infogar du en pil med dubbelt streck till vänster som ofta används i logiken.  
I kommandofönstret skriver du dlarrow.  
dubbelpil till vänster och till höger  
Med den här ikonen infogar du en pil med dubbelt streck till vänster och till höger.  
Du kan också skriva dlrarrow i kommandofönstret.  
dubbelpil till höger  
Med den här ikonen infogar du en pil med dubbelt streck till höger.  
Du kan också skriva drarrow i kommandofönstret.  
Om du vill skapa en "är mycket större än "-relation med två platshållare, skriver du <?>gg<?> eller >>.  
Med ll eller << infogar du en "är mycket mindre än "-relation i dokumentet.  
Du gör inmatningen med två platshållare enligt mönstret <?>ll<?>.  
Relationen "är definierad som" med två platshållare infogar du med hjälp av <?>def<?>.  
Ett korrespondenstecken "bild av" med två platshållare infogar du med kommandot <?>transl<?> i dokumentet.  
Kommandot <?>transr<?> infogar ett korrespondenstecken "original till" med två platshållare.  
När Du skriver in något manuellt i kommandofönstret bör Du tänka på att blankstegen är absolut nödvändiga för att Du ska åstadkomma korrekt uppbyggnad för många operatorer.  
I synnerhet gäller detta om Du arbetar med värden i stället för med platshållare, t ex om Du för relationen "är mycket större än" skulle skriva 10 gg 1 eller a gg b.  
Operatorer  
Välj den operator som du vill använda i din %PRODUCTNAME Math -formel.  
Alla tillgängliga operatorer hittar du i urvalsfönstrets nedre del.  
En motsvarande lista visas även om du öppnar snabbmeny n i fönstret Kommandon.  
Operatorer som du inte kan nå via urvalsfönstret måste du skriva in direkt i kommandofönstret.  
Alla infogningar för vilka det finns ikoner kan du givetvis även göra manuellt.  
Enbart de operatorer som listas tillsammans med en ikon kan infogas via urvalsfönstret (meny Visa - Urval) och kommandofönstrets snabbmeny.  
De olika operatorerna är:  
Limes  
Med den här ikonen infogar du tecknet för "limes av x" (gränsvärde) med en platshållare.  
Du kan också skriva lim <?> i kommandofönstret.  
Summa  
Med den här ikonen infogar du ett summatecken med en platshållare.  
I stället för att använda ikonen kan du skriva sum <?> i kommandofönstret.  
Produkt  
Med den här ikonen infogar du ett produkttecken med en platshållare.  
Du kan också skriva prod <?> i kommandofönstret.  
Koprodukt  
Med den här ikonen infogar du ett koprodukttecken med en platshållare.  
Du kan också skriva coprod <?> i kommandofönstret.  
nedre och övre gräns  
Med den här ikonen infogar du en områdesdefinition "nedre och övre gräns" för integral och summa med platshållare.  
Du kan också skriva from{ <?>} to{<?>} <?> i kommandofönstret.  
Det är bara meningsfullt att ange gränser i samband med lämpliga operatorer, jfr sum from{ <?>} to{<?>} <?>.  
Gränserna centreras över / under summatecknet.  
Integral  
Med den här ikonen infogar du en integral med en platshållare.  
Du kan också skriva int <?> i kommandofönstret.  
Dubbel integral  
Med den här ikonen infogar du en dubbel integral med en platshållare.  
Du kan också skriva iint <?> i kommandofönstret.  
Trippelintegral  
Med den här ikonen infogar du ett trippelintegraltecken med en platshållare.  
Du kan också skriva iiint <?> i kommandofönstret.  
nedre gräns  
Med den här ikonen infogar du områdesdefinitionen "nedre gräns" för integral och summa med platshållare.  
Du kan också skriva from {<?> }<?> i kommandofönstret.  
Det är bara meningsfullt att ange gränser i samband med lämpliga operatorer.  
Kurvintegral  
Med den här ikonen infogar du en kurvintegral med en platshållare.  
Du kan också skriva lint <?> i kommandofönstret.  
Dubbel kurvintegral  
Med den här ikonen infogar du en dubbel kurvintegral med en platshållare.  
I stället för att använda ikonen kan du skriva llint <?> i kommandofönstret.  
Tredubbel kurvintegral  
Med den här ikonen infogar du en tredubbel kurvintegral med en platshållare.  
Du kan också skriva lllint <?> i kommandofönstret.  
Övre gräns  
Med den här ikonen infogar du områdesdefinitionen "övre gräns" för integral och summa med platshållare.  
Du kan också skriva to {<?> }<?> i kommandofönstret.  
Det är bara meningsfullt att ange gränser i samband med lämpliga operatorer.  
Det finns ett snabbare sätt, än att skriva direkt i kommandofönstret, när Du vill förse en operator, t ex en integral, med gränser (platshållare).  
Klicka först på den önskade integralen och sedan på ikonen för gränserna.  
Limes inferior med platshållare infogar du genom att skriva liminf <?>.  
Limes superior infogar du med platshållare genom att skriva limsup <?>.  
Med oper kan du använda användardefinierade operatorer i %PRODUCTNAME Math.  
Det här alternativet är bl.a. användbart om du vill bygga in speciella tecken i en formel.  
Den här typen av operator använder du enligt följande mönster: oper %theta x.  
Den här operatorn är särskilt intressant eftersom du kan använda den för att infoga tecken som inte kommer från %PRODUCTNAME. oper kan du även använda i samband med gränser, t.ex. oper %förenar from {i=1} to n x_{i}.  
I det här exemplet finns föreningstecknet union som symbol med namnet förenar.  
Som standard är dock kommandot union inte definierat som symbol med detta namn.  
Men det går att ändra på:  
Öppna dialogrutan Symboler (menyn Verktyg - Symboler - Katalog...).  
Klicka på kommandoknappen Redigera..., varvid dialogrutan Redigera symboler öppnas.  
Välj symbolsetet special och tilldela ett lämpligt namn i kombinationsfältet Symbol, t.ex. "förenar".  
Klicka sedan på tecknet i symbolsetets visningsfält.  
Klicka först på kommandoknappen Lägg till och sedan på OK.  
Stäng dialogrutan Symboler med Stäng.  
Sedan kan du skriva tecknet i kommandofönstret enligt ovanstående mönster.  
Gränser kan även placeras på annat sätt än centrerat över / under operatorn.  
Använd de möjligheter som %PRODUCTNAME Math erbjuder för upphöjda - och nedsänkta index.  
Ange t.ex. sum_a^b c i kommandofönstret om gränserna ska justeras mot höger vid summatecknet.  
Om dina gränsdefinitioner består av längre uttryck, måste du sätta dem inom grupperingsparenteser, t.ex. sum_{ i=1}^{2*n} b.  
När du importerar formler från äldre versioner sker det automatiskt.  
Avstånden som tecknen har till varandra kan du ändra i menyerna Format - Avstånd - Kategori - Index och Format - Avstånd - Kategori - Gränser.  
Grundläggande information om index finns på ett annat ställe i hjälpen.  
När Du skriver in något manuellt i kommandofönstret bör Du tänka på att blankstegen är absolut nödvändiga för att Du ska åstadkomma korrekt uppbyggnad för många operatorer.  
Detta gäller i synnerhet om Du förser operatorerna med värden i stället för med platshållare, t ex lim a_{ n }=a.  
Funktioner  
Välj en funktion i den undre delen av fönstret.  
En lista visas om du öppnar snabbmeny n i fönstret Kommandon.  
Funktioner som inte finns i urvalsfönstret måste du skriva in direkt i kommandofönstret.  
Enbart de funktioner som listas tillsammans med en ikon kan Du infoga via urvalsfönstret (meny Visa - Urval) och kommandofönstrets snabbmeny.  
De olika funktionerna är:  
Exponentialfunktion  
Med den här ikonen infogar du en naturlig exponentialfunktion.  
I kommandofönstret kan du skriva func e^{ <?>}.  
Naturlig logaritm  
Med den här ikonen infogar du tecknet för en naturlig logaritm med platshållare.  
Om du vill infoga en sådan manuellt, skriver du ln( <?>).  
Exponentialfunktion  
Med den här ikonen infogar du en allmän exponentialfunktion med platshållare.  
Samma resultat får du om du skriver exp( <?>) i kommandofönstret.  
Logaritm  
Med den här ikonen infogar du tecknet för en logaritm.  
Samma tecken infogas om du skriver log( <?>) manuellt.  
Potens  
Med den här ikonen infogar du en variabel med exponent till höger.  
Du kan också skriva <?>^{ <?>} i kommandofönstret. ^ -tecknet kan du ersätta med rsup eller sup.  
Sinus  
Med den här ikonen infogar du ett sinustecken med en platshållare.  
Du kan också skriva sin( <?>) i kommandofönstret.  
Cosinus  
Med den här ikonen infogar du ett cosinustecken med en platshållare.  
Du kan också skriva cos( <?>) i kommandofönstret.  
Tangens  
Med den här ikonen infogar du ett tangenstecken med en platshållare.  
Du kan också skriva tan (<?>) i kommandofönstret.  
Cotangens  
Med den här ikonen infogar du ett cotangenstecken med en platshållare.  
Du kan också skriva cot( <?>) i kommandofönstret.  
Hyperbolisk sinus  
Med den här ikonen infogar du ett tecken för hyperbolisk sinus med en platshållare.  
Du kan också skriva sinh( <?>) i kommandofönstret.  
Kvadratrot  
Med den här ikonen infogar du en kvadratrot med platshållare.  
Vid direkt inmatning i kommandofönstret skriver du sqrt <?>.  
Hyperbolisk cosinus  
Med den här ikonen infogar du ett tecken för hyperbolisk cosinus med en platshållare.  
Du kan också skriva cosh( <?>) i kommandofönstret.  
Hyperbolisk tangens  
Med den här ikonen infogar du ett tecken för hyperbolisk tangens med en platshållare.  
Du kan också skriva tanh( <?>) i kommandofönstret.  
Hyperbolisk cotangens  
Med den här ikonen infogar du ett tecken för hyperbolisk cotangens med en platshållare.  
Du kan också skriva coth( <?>) i kommandofönstret.  
N-te roten  
Med den här ikonen infogar du tecknet för n-te rot ur x med två platshållare.  
Samma resultat får du om du skriver nroot n x i kommandofönstret.  
Arcussinus  
Med den här ikonen infogar du ett arcussinustecken med en platshållare.  
Du kan också skriva arcsin( <?>) i kommandofönstret.  
Arcuscosinus  
Med den här ikonen infogar du ett arcuscosinustecken med en platshållare.  
Du kan också skriva arccos( <?>) i kommandofönstret.  
Arcustangens  
Med den här ikonen infogar Du tecknet för arcustangens med en platshållare.  
Du kan också skriva arctan( <?>) i kommandofönstret.  
Arcuscotangens  
Med den här ikonen infogar du tecknet för arcuscotangens med en platshållare.  
Du kan också skriva arccot( <?>) i kommandofönstret.  
Absolutvärde  
Med den här ikonen infogar du ett absolutvärde med platshållare.  
I stället för att använda ikonen kan du skriva abs <?> direkt i kommandofönstret.  
Area sinus hyperbolicus  
Med den här ikonen infogar Du tecknet för area sinus hyperbolicus med en platshållare.  
Du kan också skriva arsinh( <?>) i kommandofönstret.  
Area cosinus hyperbolicus  
Med den här ikonen infogar du tecknet för area cosinus hyperbolicus med en platshållare.  
Du kan också skriva arcosh( <?>) i kommandofönstret.  
Area tangens hyperbolicus  
Med den här ikonen infogar du tecknet för area tangens hyperbolicus med en platshållare.  
I stället för att använda ikonen kan du skriva artanh( <?>) i kommandofönstret.  
Area cotangens hyperbolicus  
Med den här ikonen infogar du tecknet för area cotangens hyperbolicus med en platshållare.  
I stället för att använda ikonen kan du skriva arcoth( <?>) i kommandofönstret.  
Fakultet  
Med den här ikonen infogar du ett fakultetstecken med platshållare.  
I stället för att använda ikonen kan du skriva fact <?> i kommandofönstret.  
Du kan även förse en funktion med index eller exponent.  
Testa själv genom att mata in följande i kommandofönstret: sin^2x+cos^2x=1.  
Även funktionen func f_x def{ partial func f}over{partial x} är ett bra exempel på detta.  
När du matar in funktioner manuellt i kommandofönstret bör du tänka på att mellanslag är absolut nödvändiga för vissa funktioner. (t.ex. abs 5=5; abs -3=3)  
Parenteser  
Välj den parentes som du vill använda i din %PRODUCTNAME Math -formel.  
Parenteserna som är tillgängliga i urvalsfönstret finns i fönstrets nedre del.  
En motsvarande lista visas även om du öppnar snabbmeny n i fönstret Kommandon.  
Parenteser som du inte kan nå via urvalsfönstret måste du skriva in direkt i kommandofönstret.  
Du kan givetvis göra alla infogningar manuellt, även om det finns ikoner till dem.  
Det är bara parenteser med en ikon som du kan infoga via urvalsfönstret (menyn Visa - Urval) snabbmenyn i kommandofönstret.  
De olika parenteserna är:  
Parenteser  
Med den här ikonen infogar du en platshållare omgiven av normala runda parenteser.  
Du kan också skriva (<?>) direkt i kommandofönstret.  
Hakparenteser  
Med den här ikonen infogar du en platshållare omgiven av hakparenteser.  
Du kan också skriva [<?>] direkt i kommandofönstret.  
Dubbla hakparenteser  
Med den här ikonen infogar du en platshållare omgiven av dubbla hakparenteser.  
Du kan också skriva ldbracket <?> rdbracket direkt i kommandofönstret.  
Klammerparenteser  
Med den här ikonen infogar du en platshållare omgiven av klammerparenteser.  
I stället för att använda ikonen kan du skriva lbrace<?>rbrace direkt i kommandofönstret.  
Enkla linjer  
Med den här ikonen infogar du en platshållare omgiven av enkla linjer.  
I stället för att använda ikonen kan du skriva lline <?> rline direkt i kommandofönstret.  
Dubbla linjer  
Med den här ikonen infogar du en platshållare omgiven av dubbla linjer.  
I stället för att använda ikonen kan du skriva ldline<?>rdline direkt i kommandofönstret.  
Vinkelparenteser  
Med den här ikonen infogar du en platshållare omgiven av vinkelparenteser.  
I stället för att använda ikonen kan du skriva langle<?> rangle direkt i kommandofönstret.  
Operatorparenteser  
Med den här ikonen infogar du operatorparenteser, d.v.s. vinkelparenteser med platshållare.  
I stället för att använda ikonen kan du skriva langle <?> mline <?> rangle i kommandofönstret.  
Grupperingsparenteser  
Med den här ikonen infogar du grupperingsparenteser.  
I stället för att använda ikonen kan du skriva {<?>} direkt i kommandofönstret.  
Parenteser (skalbara)  
Med den här ikonen infogar du runda vänster och höger parenteser med platshållare.  
I stället för att använda ikonen kan du skriva left( <?> right) i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Vänster och höger hakparentes  
Med den här ikonen infogar du hakparenteser med platshållare.  
I stället för att använda ikonen kan du skriva left[ <?> right] direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Dubbla hakparenteser (skalbara)  
Med den här ikonen infogar du dubbla hakparenteser med platshållare.  
I stället för att använda ikonen kan du skriva left ldbracket <?> right rdbracket direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Vänster och höger klammerparentes  
Med den här ikonen infogar du skalbara klammerparenteser med platshållare.  
I stället för att använda ikonen kan du skriva left lbrace <?> right rbrace direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Enkla linjer (skalbara)  
Med den här ikonen infogar du skalbara vänster - och högerlinjer med platshållare.  
I stället för att använda ikonen kan du skriva left lline <?> right rline direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Med "a" menas platshållaren som du tilldelar respektive formatering.  
Givetvis kan du ersätta den med valfria tecken.  
Med den här ikonen infogar du en platshållare omgiven av dubbla linjer.  
I stället för att använda ikonen kan du skriva left ldline<?> right rdline direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Vinkelparenteser (skalbara)  
Med den här ikonen infogar du skalbara vinkelparenteser med platshållare.  
I stället för att använda ikonen kan du skriva left langle <?> right rangle direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Operatorparenteser (skalbara)  
Med den här ikonen infogar du operatorparenteser (skalbara), d.v.s. skalbara vinkelparenteser med platshållare.  
I stället för att använda ikonen kan du skriva left langle <?> mline <?> right rangle direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Klammerparentes uppe (skalbar)  
Med den här ikonen infogar du en skalbar horisontell klammerparentes uppe med platshållare.  
I stället för att använda ikonen kan du skriva <?> overbrace <?> direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Klammerparentes nere (skalbar)  
Med den här ikonen infogar du en skalbar horisontell klammerparentes nere med platshållare.  
I stället för att använda ikonen kan du skriva <?> underbrace <?> direkt i kommandofönstret.  
Parentesernas storlek anpassas automatiskt.  
Vid direkt inmatning i kommandofönstret infogar du vänster - och högerlinjer med kanter nedtill och en platshållare mellan dem genom att skriva lfloor<?>rfloor.  
Men du kan även skriva in detta utan platshållartecken.  
Vid direkt inmatning i kommandofönstret infogar du vänster - och högerlinjer med kanter upptill och en platshållare mellan dem genom att skriva lceil<?>rceil.  
Du kan även skriva in detta utan platshållartecken.  
Linjerna anpassas automatiskt till teckenstorleken.  
Du kan även skriva in detta utan platshållar-tecken.  
Linjerna anpassas automatiskt till teckenstorleken.  
Du kan även skriva in detta utan platshållartecken.  
Storleken på parenteser anpassas automatiskt om du skriver left och right framför parenteserna, t.ex. left( a over b right).  
Du kan göra inställningar av storleksanpassningen om du väljer Format - Avstånd... - Kategori - Parenteser.  
I fältet Vänster / höger överstorlek anger du t.ex. 5 procent som storlek.  
Sedan markerar du fältet Skala alla parenteser och ställer in 0 procent i det tillhörande rotationsfältet Överstorlek.  
Följande exempel demonstrerar resultatet av en inställningen av den här typen: left (left (left ((((a over b))) right) right) right).  
Samtliga parenteser går även att använda utan grupperingsfunktion, d.v.s. enskilt.  
Då måste du placera det omvända snedstrecket\ (backslash) framför respektive kommando.  
Om du t.ex. skriver\ [, så visas den vänstra hakparentesen utan dess högra motsvarighet.  
Med snedstrecket kan du alltså även byta plats på parenteser.  
Om du skriver\]\ [placeras hakparenteserna med baksidorna mot varandra.  
Detta har du bl.a. nytta av om du vill bygga upp intervaller.  
Prova följande exempel för ett öppet intervall:\] a;b\[=lbrace x \lline a<x<b rbrace. (Du kan kopiera formeln här och klistra in den i kommandofönstret.) Men det är bara de icke-skalbara parenteserna som kan användas var för sig.  
Om du vill ändra storleken, måste du använda kommandot size enligt mönstret size 50\ [.  
När du skriver in något direkt i kommandofönstret bör du tänka på att mellanslag är absolut nödvändiga i vissa parenteser för den korrekta uppbyggnaden, t.ex. left ldline<?> right rdline.  
Mer information om formatering i %PRODUCTNAME Math får du om du klickar på den här hyperlänken.  
Med hjälp av informationen om Index och exponenter och Skalning kan du ge dina dokument en optimal utformning.  
Det finns även mer information om Parenteser och grupperingar.  
Attribut  
Tilldela tecknen i din %PRODUCTNAME Math -formel olika attribut.  
I urvalsfönstrets nedre del visas de olika attributen.  
Du kan även visa motsvarande lista genom att öppna snabbmeny n i fönstret Kommandon.  
Attribut som du inte kan nå via urvalsfönstret måste du skriva in direkt i kommandofönstret.  
Du kan givetvis även göra alla infogningar manuellt, även dem för vilka det finns ikoner.  
Det är bara de attribut som listas tillsammans med en ikon som du kan infoga via urvalsfönstret (menyn Visa - Urval) och kommandofönstrets snabbmeny.  
Med "a" menas en platshållare som du tilldelar respektive attribut.  
Givetvis kan du ersätta den med valfria tecken.  
De olika attributen är:  
Accent åt höger  
Med den här ikonen infogar du en platshållare med en accent åt höger (akut).  
I stället för att använda ikonen kan du skriva acute<?> direkt i kommandofönstret.  
Accent åt vänster  
Med den här ikonen infogar du en platshållare med en accent åt vänster (grav).  
I stället för att använda ikonen kan du skriva grave<?> direkt i kommandofönstret.  
Omvänd cirkumflex  
Med den här ikonen infogar du en platshållare med en omvänd cirkumflex ovanför.  
I stället för att använda ikonen kan du skriva check<?> direkt i kommandofönstret.  
Breve  
Med den här ikonen infogar du en platshållare med breve (korttecken).  
I stället för att använda ikonen kan du skriva breve<?> direkt i kommandofönstret.  
Cirkel  
Med den här ikonen infogar du en platshållare med en cirkel ovanför.  
I stället för att använda ikonen kan du skriva circle <?> direkt i kommandofönstret.  
Vektorpil  
Med den här ikonen infogar du en platshållare med en vektorpil.  
I stället för att använda ikonen kan du skriva vec<?> direkt i kommandofönstret.  
Tilde  
Med den här ikonen infogar du en platshållare med en tilde.  
I stället för att använda ikonen kan du skriva tilde<?> direkt i kommandofönstret.  
Cirkumflex  
Med den här ikonen infogar du en platshållare med en cirkumflex (ett "tak") ovanför.  
I stället för att använda ikonen kan du skriva hat<?> direkt i kommandofönstret.  
Linje över  
Med den här ikonen infogar du en platshållare med en linje ovanför.  
I stället för att använda ikonen kan du skriva bar<?> direkt i kommandofönstret.  
Det här attributet påverkar bara ett tecken.  
Punkt  
Med den här ikonen infogar du en platshållare med en punkt ovanför.  
I stället för att använda ikonen kan du skriva dot<?> i kommandofönstret.  
Bred vektorpil  
Med den här ikonen infogar du en bred vektorpil med platshållare.  
I stället för att använda ikonen kan du skriva widevec direkt i kommandofönstret.  
Bred tilde  
Med den här ikonen infogar du en bred tilde med platshållare.  
Du kan också skriva widetilde direkt i kommandofönstret.  
Bred cirkumflex  
Med den här ikonen infogar du en bred cirkumflex med en platshållare.  
I stället för att använda ikonen kan du skriva widehat direkt i kommandofönstret.  
Dubbel punkt  
Med den här ikonen infogar du en platshållare med två punkter ovanför.  
I stället för att använda ikonen kan du skriva ddot<?> direkt i kommandofönstret.  
Linje över  
Med den här ikonen infogar du en platshållare med en upphöjd linje ovanför.  
I stället för att använda ikonen kan du skriva overline<?> direkt i kommandofönstret.  
Linjens längd anpassar sig till antalet tecken.  
Linje under  
Med den här ikonen infogar du en platshållare med en nedsänkt linje nedanför.  
I stället för att använda ikonen kan du skriva underline<?> direkt i kommandofönstret.  
Linje genom  
Med den här ikonen infogar du en platshållare med en linje genom.  
I stället för att använda ikonen kan du skriva overstrike<?> direkt i kommandofönstret.  
Tredubbel punkt  
Med den här ikonen infogar du en platshållare med tre punkter ovanför.  
I stället för att använda ikonen kan du skriva dddot<?> direkt i kommandofönstret.  
Transparent  
Med den här ikonen infogar du en platshållare med ett transparent tecken som upptar samma utrymme som a men som inte visas.  
I stället för att använda ikonen kan du skriva phantom <?> direkt i kommandofönstret.  
Fetstil  
Med den här ikonen infogar du en platshållare med formatet fet.  
I stället för att använda ikonen kan du skriva bold<?> i kommandofönstret.  
Kursivt teckensnitt  
Med den här ikonen infogar du en platshållare med formatet kursiv.  
I stället för att använda ikonen kan du skriva ital <?> eller italic direkt i kommandofönstret.  
Ändra storlek  
Med den här ikonen infogar du kommandot som ändrar teckenstorlek med två platshållare.  
Den första platshållaren innehåller teckenstorleken, t.ex. 12, den andra innehåller texten.  
Glöm inte att foga in blanksteg mellan värdena.  
I stället för att använda ikonen kan du skriva size<?> <?> direkt i kommandofönstret.  
Det är meningslöst att använda kommandot size fristående.  
Ändra teckensnitt  
Med den här ikonen infogar du kommandot som ändrar teckensnitt med två platshållare.  
För den första platshållaren använder du ett av namnen för användarteckensnitten Serif, Sans eller Fixed.  
Den andra platshållaren innehåller den formaterade texten.  
I ställer för att använda ikonen kan du skriva font<?><?> direkt i kommandofönstret.  
Fristående, d.v.s. utan tecken som ska formateras, är kommandot font meningslöst.  
Om du vill visa tecken i färg i en formel använder du kommandot color.  
Du måste ange kommandot tillsammans med någon av de tillgängliga färgerna white, black, cyan, magenta, red, blue, green eller yellow, följt av ett tecken eller en sammanhörande teckenföljd.  
Följande exempel belyser detta: color green size 20 a.  
Lägg märke till att två attribut (färg och storlek) används för bokstaven a.  
Om delar av formeln har formaterats feta eller kursiva av programmet och du vill ta bort dessa attribut, kan du använda kommandona nbold och nitalic.  
Ska t.ex. tecknet x i formeln 5 x + 3=28 inte längre vara kursivt, måste du infoga nitalic framför x, d.v.s. du måste skriva 5 nitalic x + 3=28.  
Attributen "acute", "bar", "breve", "check", "circle", "dot", "ddot", "dddot", "grave", "hat", "tilde" och "vec "har fasta storlekar.  
De blir inte bredare respektive längre om de står över en lång symbol.  
När Du vill ändra storlek kan Du använda size n, +n, -n, *n och / n, varvid n fungerar som platshållare.  
Formerna med "förtecken" är särskilt lämpliga när Du ska göra eventuella ändringar av basstorleken.  
Du kan kopiera och infoga dem på annat ställe utan att deras utseende ändras.  
Med size +n och size -n ändrar Du storleken i punkter (pt, points).  
Procentuella ändringar åstadkommer Du med size *n och size / n, varvid snedstrecket får proportionella förhållanden.  
Om Du t ex vill förstora ett tecken med 17%, måste Du skriva size *1.17.  
När Du skriver in något manuellt i kommandofönstret bör Du tänka på att blankstegen ibland är absolut nödvändiga för att kommandot ska byggas upp korrekt.  
I synnerhet gäller detta om Du förser Dina attribut med värden i stället för med platshållare, t ex font sans 20.  
Du får mer information om formatering i %PRODUCTNAME Math om du klickar på den här hyperlänken.  
Värdefull information om attribut, index och exponenter samt skalning hjälper dig att utforma dina dokument optimalt.  
Formateringar  
Här hittar du många alternativ med vars hjälp du kan justera tecknen i %PRODUCTNAME Math -formeln optimalt.  
I urvalsfönstrets nedre del visas de olika justeringsmöjligheterna.  
Du kan även visa en lista med samma funktioner om du öppnar snabbmeny n i fönstret Kommandon.  
Det är bara formateringarna som listas tillsammans med en ikon som du kan infoga via urvalsfönstret (menyn Visa - Urval) och snabbmenyn i kommandofönstret.  
Med "a" menas alltid den platshållare i formeln som Du vill tilldela den aktuella formateringen.  
Du kan skriva ett valfritt tecken.  
De olika formateringarna är:  
Exponent till vänster  
Med den här ikonen infogar du en variabel med exponent till vänster och en platshållare.  
I stället för att använda ikonen kan du skriva <?>lsup{ <?>} i kommandofönstret.  
Exponent uppe  
Med den här ikonen infogar du en exponent direkt över en variabel.  
I stället för att använda ikonen kan du skriva <?>csup <?> direkt i kommandofönstret.  
Exponent till höger  
Med den här ikonen infogar du en variabel med exponent till höger.  
I stället för att använda ikonen kan du skriva <?>^{ <?>} i kommandofönstret. ^ -tecknet kan du ersätta med rsup eller sup.  
Vertikal placering (två element)  
Med den här ikonen infogar du ett binom med två platshållare.  
I stället för att använda ikonen kan du skriva binom<?><?> i kommandofönstret.  
Börja ny rad  
Med den här ikonen infogar du en ny rad i dokumentet.  
I stället för att använda ikonen kan du skriva newline direkt i kommandofönstret.  
Index till vänster  
Med den här ikonen infogar du en variabel med index till vänster och en platshållare.  
I stället för att använda ikonen kan du skriva <?>lsub{ <?>} direkt i kommandofönstret.  
Index nere  
Med den här ikonen infogar du ett index direkt under en variabel.  
I stället för att använda ikonen kan du skriva csub direkt i kommandofönstret.  
Du gör inmatningen enligt mönstret <?>csub <?>.  
Index till höger  
Med den här ikonen infogar du en variabel med index.  
I stället för att använda ikonen kan du skriva <?>_{ <?>} direkt i kommandofönstret.  
Du kan ersätta det nedsänkta strecket med rsub eller sub.  
Vertikal placering (tre element)  
Med den här ikonen infogar du en stack med tre platshållare.  
I stället för att använda ikonen kan du skriva stack {<?>#<?>#<?>} direkt i kommandofönstret.  
Litet mellanrum  
Med den här ikonen infogar du ett litet mellanslag med platshållare.  
I stället för att använda ikonen kan du skriva tecknet ` direkt i kommandofönstret.  
Men det är bara meningsfullt om det står till vänster eller höger om en symbol, en variabel, ett tal eller ett fullständigt kommando.  
Vänsterjustera  
Med den här ikonen infogar du kommandot för vänsterjustering av "a" med en platshållare.  
I stället för att använda ikonen kan du skriva alignl<?> direkt i kommandofönstret.  
Justera centrerat (horisontellt)  
Med den här ikonen infogar du kommandot för en horisontell centrering av "a" med en platshållare.  
I stället för att använda ikonen kan du skriva alignc<?> direkt i kommandofönstret.  
Högerjustera  
Med den här ikonen infogar du kommandot för högerjustering av "a" med en platshållare.  
I stället för att använda ikonen kan du skriva alignr<?> direkt i kommandofönstret.  
Matrisplacering  
Med den här ikonen infogar du en matris med fyra platshållare.  
I stället för att använda ikonen kan du skriva matrix {<?>#<?>##<?>#<?>#} direkt i kommandofönstret.  
Det första tecknet anger radnumret och det andra tecknet kolumnnumret där elementet står.  
Du kan utöka matrisen i kommandofönstret genom att infoga fler tecken.  
Mellanrum  
Med den här ikonen infogar du ett mellanslag med platshållare.  
I stället för att använda ikonen kan du skriva en tilde ~ direkt i kommandofönstret.  
Men det är bara meningsfullt om det finns en symbol, en variabel, ett tal eller ett fullständigt kommando till vänster eller höger om tilden.  
Justering med kommandona alignl, alignc och alignr är särskilt effektiv om du  
justerar täljare och nämnare, t ex {alignl a}over{b+c},  
bygger upp binom eller stackar, t ex binom{ 2*n}{alignr k},  
justerar elementen i en matris, t ex matrix{ alignr a#b+2##c+1 / 3#alignl d} eller  
börjar en ny rad, t ex a+b-c newline alignr x / y.  
När Du använder align-instruktioner måste Du tänka på att dessa  
bara får stå i början på uttryck, och dessutom bara en gång.  
Du kan alltså inte skriva a+alignr b. medan däremot a+b alignr c  
påverkar varandra, vilket leder till att a justeras mot höger när Du anger {alignl{alignr a}}over{b+c}.  
Om en rad eller ett uttryck börjar med text, så vänsterjusteras raden / stycket som standard.  
Med motsvarande align-kommandon kan Du givetvis utföra en avvikande formatering, jfr stack{ a+b-c*d#a-b+c#"text"} med stack{a+b-c*d#alignl a-b+c#alignr "text"}.  
Text måste alltid inneslutas av citattecken (dock inte typografiska).  
Du kan utnyttja tomma grupper eller strängar vid justering på ett intressant sätt.  
Placera en tom sträng, dvs de citattecken "" som innesluter varje text, framför den formeldel som Du vill justera mot vänster.  
Formler centreras som standard men Du kan justera dem mot vänster utan att använda menyn Format - Justering, jfr "Ett exempel" newline a+b newline ""c-d.  
Du kan göra likadant med tomma grupper, jfr b+b+b+b+{ }"Detta är ytterligare ett exempel "newline a+a+a+a+a+a.  
Här kommer texten, under förutsättning att standardinställningen inte har ändrats, också att centreras.  
När Du skriver in något manuellt i kommandofönstret bör Du tänka på att blankstegen i vissa formateringar är absolut nödvändiga för att kommandot ska byggas upp korrekt.  
Detta gäller i synnerhet om Du anger värden i stället för platshållare, t ex a lsup{ 3}.  
Du får mer information om formatering i %PRODUCTNAME Math om du klickar på den här hyperlänken.  
Med hjälp av mer information om Index och exponenter och Skalning kan du ge dina dokument en optimal utformning.  
Mängdoperationer  
Tilldela tecknen i din %PRODUCTNAME Math -formel olika mängdoperatorer.  
De olika operatorerna visas i nedre delen av urvalsfönstret.  
Du kan även visa en lista med samma funktioner genom att öppna snabbmeny n i fönstret Kommandon.  
Alla operatorer som inte finns med i urvalsfönstret måste du ange direkt i kommandofönstret.  
Du kan göra alla infogningar direkt, även dem för vilka det finns ikoner.  
När du klickar på ikonen Mängdoperationer visas fler symboler.  
Du kan infoga dessa symboler i formeln i kommandofönstret genom att klicka på dem.  
De olika mängdoperationerna är:  
finns i  
Med den här ikonen infogar du mängdoperatorn "finns i" med två platshållare.  
I stället för att använda ikonen kan du skriva <?> in <?> i kommandofönstret.  
finns inte i  
Med den här ikonen infogar du mängdoperatorn "finns inte i" med två platshållare.  
I stället för att använda ikonen kan du skriva <?> notin <?> direkt i kommandofönstret.  
innehåller  
Med den här ikonen infogar du mängdoperatorn innehåller med två platshållare.  
Om du använder kommandona owns eller ni, måste du ange dem enligt mönstret <?>ni<?>.  
Tom mängd  
Med den här ikonen infogar du en tom mängd.  
I stället för att använda ikonen kan du skriva emptyset direkt i kommandofönstret.  
Genomsnitt  
Med den här ikonen infogar du två platshållare med mängdoperatorn genomsnitt av mängder.  
I stället för att använda ikonen kan du skriva <?>intersection<?> direkt i kommandofönstret.  
Union  
Med den här ikonen infogar du mängdoperatorn "union av mängder" med två platshållare i dokumentet.  
I stället för att använda ikonen kan du skriva <?>union<?> direkt i kommandofönstret.  
Differens  
Med den här ikonen infogar du mängdoperatorn "differens av mängder" i dokumentet.  
Du måste ange dem enligt mönstret <?>setminus<?>.  
Kvotmängd  
Med den här ikonen infogar du / -tecknet för uppbyggnad av en kvotmängd med två platshållare.  
I stället för att använda ikonen kan du skriva <?>slash<?> direkt i kommandofönstret.  
Alef  
Med den här ikonen infogar du ett kardinaltal.  
I stället för att använda ikonen kan du skriva aleph i kommandofönstret.  
Delmängd  
Med den här ikonen infogar du mängdoperatorn "är delmängd av".  
I stället för att använda ikonen kan du skriva <?>subset<?> direkt i kommandofönstret.  
Delmängd eller lika  
Med den här ikonen infogar du mängdoperatorn "delmängd eller lika" med två platshållare.  
I stället för att använda ikonen kan du skriva <?>subseteq<?> direkt i kommandofönstret.  
Grundmängd  
Med den här ikonen infogar du mängdoperatorn "är grundmängd av" och två platshållare.  
I stället för att använda ikonen kan du skriva <?>supset<?> direkt i kommandofönstret.  
Grundmängd eller lika  
Med den här ikonen infogar du mängdoperatorn "är grundmängd eller lika" med två platshållare.  
I stället för att använda ikonen kan du skriva <?>supseteq<?> direkt i kommandofönstret.  
Inte delmängd  
Med den här ikonen infogar du mängdoperatorn "inte delmängd" med två platshållare.  
I stället för att använda ikonen kan du skriva <?>nsubset<?> direkt i kommandofönstret.  
Inte delmängd eller lika  
Med den här ikonen infogar du mängdoperatorn "inte delmängd eller lika" med två platshållare.  
I stället för att använda ikonen kan du skriva <?>nsubseteq<?> direkt i kommandofönstret.  
Inte grundmängd  
Med den här ikonen infogar du mängdoperatorn "inte grundmängd" med två platshållare.  
I stället för att använda ikonen kan du skriva <?>nsupset<?> direkt i kommandofönstret.  
Inte grundmängd eller lika  
Med den här ikonen infogar du mängdoperatorn "inte grundmängd eller lika" med två platshållare.  
I stället för att använda ikonen kan du skriva <?>nsupseteq<?> direkt i kommandofönstret.  
Mängd naturliga tal  
Med den här ikonen infogar du ett tecken för "mängd naturliga tal".  
I stället för att använda ikonen kan du skriva setn direkt i kommandofönstret.  
Heltalsmängd  
Med den här ikonen infogar du ett tecken för heltalsmängd.  
I stället för att använda ikonen kan du skriva setz direkt i kommandofönstret.  
Mängd rationella tal  
Med den här ikonen infogar du ett tecken för Mängd rationella tal.  
I stället för att använda ikonen kan du skriva setq direkt i kommandofönstret.  
Mängd reella tal  
Med den här ikonen infogar du ett tecken för mängd reella tal.  
I stället för att använda ikonen kan du skriva setr direkt i kommandofönstret.  
Mängd komplexa tal  
Med den här ikonen infogar du ett tecken för mängd komplexa tal.  
I stället för att använda ikonen kan du skriva setc direkt i kommandofönstret.  
När Du skriver in något manuellt i kommandofönstret bör Du tänka på att blankstegen är absolut nödvändiga för att Du ska åstadkomma korrekt uppbyggnad för många operatorer.  
Detta gäller i synnerhet om Du arbetar med värden i stället för med platshållare, t ex om Du i stället för mängdoperatorn delmängd skriver A subset B.  
Exempel  
Här får du några exempelformler för det dagliga arbetet med %PRODUCTNAME Math.  
Symbol med index  
Här hittar du ett exempel på hur du skapar symboler med index med %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax:  
D_{ mn}^ {size / 2 LEFT(3 OVER 2 RIGHT)}  
Symbol med index  
Här hittar du ett andra exempel på hur du skapar symboler med index med %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax: %SIGMA_g^{ {}+{} }lsup 3  
Symbol med index  
Här hittar du ett tredje exempel på hur du skapar symboler med index med %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax: %PHI^{ i_1 i_2 dotsaxis i_n}_{k_1 k_2 dotsaxis k_n}  
Matris med olika teckenstorlekar  
Här hittar du ett exempel på hur du skapar en matris med olika teckenstorlekar i %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax: func G^{ (%alpha "," %beta)}_ {x_m x_n} = left [matrix {arctan(%alpha) # arctan(%beta) ## x_m + x_n # x_m - x_n }right]  
Matris  
Här hittar du ett exempel på hur du skapar en matris med %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax: font sans bold size *1,5 A =left[ matrix{A_11#A_12#dotsaxis#A_{1n}##A_21#{} #{}#A_{2n}##dotsvert#{}#{}#dotsvert##A_{n1}#A_{n2}#dotsaxis#A_nn}right]  
Matris med fetstil  
Här hittar du ett exempel på hur du skapar en matris med fetstil i %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax: bold {f(x", "y) = left [stack {x + y over z + left lbrace matrix {2 # 3 # 4 ## 4 # 5 # 6 ## 6 # 7 # 8} right rbrace # {y + sin (x)} over %alpha # z + y over g} right]}  
Funktion  
Här hittar du ett exempel på hur du skapar funktioner med %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax: func f( x" ,"y)={x sin x~ tan y} over {cos x}  
Kvadratrot  
Här hittar du ett exempel på hur du skapar en kvadratrot med %PRODUCTNAME Math.  
Om du vill överta exemplets syntax för ditt arbete, kan du kopiera den till fönstret Kommandon via urklippet.  
Syntax: %LAMBDA_{ deg" ,"t}=1 + %alpha_deg SQRT {M_t over M_{(t=0)}-1}~". "  
Olika teckensnitt och teckenstorlekar  
Här hittar du ett exempel på hur du använder olika teckensnitt och teckenstorlekar med %PRODUCTNAME Math.  
Syntax: f( t)=int from size*1.5 0 to 1 left[g(t')+sum from i=1 to N h_i(t')right]  
Attribut  
Här hittar du ett exempel på hur du använder olika attribut i en formel med %PRODUCTNAME Math.  
Syntax: %rho( font sans bold q" ,"%omega) = int func e^{i %omega t}%rho(font sans bold q" ,"t)"d "t  
Parenteser och grupperingar  
Citattecknen i exemplen används bara för att framhäva delar av texten och innehållsligt hör de inte till exemplen och kommandona.  
När du skriver exempel i kommandofönstret manuellt bör du tänka på att du ofta måste använda blanksteg för ge exemplen korrekt uppbyggnad.  
De viktigaste parenteserna är klammerparenteserna "{}" med vilka du kan gruppera flera uttryck / symboler till ett nytt uttryck.  
Exemplet "{a + b}over{c + d} - e" illustrerar detta.  
Parenteserna visas inte i formeldokumentet och behöver inte heller något som helst utrymme.  
Klammerparenteser har hittills infogats via urvalsfönstret eller direkt i kommandofönstret på följande sätt: "left lbrace <?> right rbrace".  
Nu kan Du även infoga en vänster och en höger klammerparentes med "lbrace" och "rbrace ", och detta med eller utan platshållare.  
Du tillgång till sammanlagt åtta (8) olika parentestyper!  
Parentestyperna "ceil" - och "floor" används ofta inom informatiken för att avrunda argument uppåt eller nedåt till närmaste heltal: "lceil -3.7 rceil = -3 "eller "lfloor -3.7 rfloor = -4".  
Vinkelparenteser med ett lodrätt streck mellan dem är rätt vanliga inom fysiken: "langle a mline b rangle" eller "langle a mline b mline c over d mline e rangle ".  
De lodräta streckens höjd och placering motsvarar alltid exakt de omgivande parenteserna.  
Alla parenteser får bara förekomma som enhetliga par.  
Parenteserna har några gemensamma drag:  
Alla parentestyper har en grupperande funktion, likt den som beskrivs för "{}" - parenteserna.  
Du kan använda alla parentestyper, dvs även de synliga, för att definiera tomma grupper.  
Det inneslutna uttrycket får alltså vara tomt.  
Ytterligare en gemensam egenskap för alla dessa parenteser är det att de inte anpassar sin storlek till det inneslutna uttrycket, vilket gäller åt båda håll.  
Om Du t ex vill visa "(a over b)" med en parentesstorlek som anpassats till a och b, så måste Du infoga "left "och "right".  
Genom att ange "left(a over b right)" får Du lämpliga storleksförhållanden.  
Samma sak gäller för de olika inmatningssätten, alltså även för de motsvarande resultaten för "(size 3{a over b})" och "left(size 3{a over b}right) ".  
Om parenteserna själva är en del av det uttryck vars storlek ändras, så berörs även de av storleksändringen: "size 3(a over b)" och "size 12(a over b) ".  
Givetvis ändrar detta inte någonting på storleksförhållandet mellan parentesen och det inneslutna uttrycket.  
Eftersom "left" och "right "säkerställer en entydig tilldelning av parenteserna till varandra, kan Du använda varje enskild parentes som argument för dessa båda, även för höger parentes på vänster sida och omvänt.  
I stället för en parentes kan det även stå "none", vilket betyder att det inte visas någon parentes på detta ställe och att det inte heller reserveras utrymme för någon parentes.  
På så vis kan Du t ex bilda följande uttryck:  
left lbrace x right none  
left [x right)  
left] x right [  
left rangle x right lfloor  
De fungerar även grupperande och får innesluta det tomma uttrycket.  
En kombination av parenteser som inte hör till varandra, samt parenteser på bara en sida och positionsbyte av höger och vänster parentes förekommer ofta.  
Ett exempel från matematiken, som dock inte kan skrivas in så, förtydligar detta:  
[2, 3) - intervall som är öppet till höger  
Men parenteserna har då inte någon fast storlek eftersom de anpassar sig till argumentet.  
Därför går det nu att visa enskilda parenteser med fast storlek genom att man sätter ett omvänt snedstreck "\" (backslash) framför de vanliga parenteserna.  
Dessa parenteser uppför sig sedan som vilken symbol som helst och har inte längre några parentesspecifika funktioner, dvs de fungerar inte grupperande och de justeras som andra symboler, jfr "size *2 \langle x \rangle" och "size *2 langle x rangle ".  
En fullständig översikt ser därför ut som följer:  
\{ eller \lbrace,\} eller \rbrace  
\(,\)  
\[,\]  
\langle, \rangle  
\lceil, \rceil  
\lfloor, \rfloor  
\lline, \rline  
\ldline, \rdline  
Därmed kan Du bygga upp sådana intervall som det ovanstående utan problem i %PRODUCTNAME Math: \[ 2", "3\) eller "\]2", "3\ [(Observera:  
Dessa citattecken hör till inmatningen.)  
Se till att du använder de citattecken som du tar fram med Skift+2 och inte de typografiska.  
Av princip bör skiljetecken (som kommatecknet i det här fallet) alltid sättas som text, även blanksteg kan ofta vara lämpliga.  
Du kan visserligen även använda "\[2,~3\)", men ovanstående möjlighet är att föredra.  
Beteckningen "fast storlek" betyder i det ovanstående alltid att parentesernas storlek bara är beroende av den använda teckenstorleken.  
Att kapsla grupperingar är relativt oproblematiskt.  
För hat "{a + b}" visas "hat", dvs circumflex (^), mitt över "{a + b} ".  
Även "color red lceil a rceil" och "grave hat langle x * y rangle "fungerar som förväntat.  
Det senare ger ett liknande resultat som "grave {hat langle x * y rangle}".  
Detta är inte överraskande, eftersom dessa attribut inte konkurrerar med varandra, utan kan kombineras.  
Något annorlunda förhåller det sig däremot med attributen, som konkurrerar med varandra eller som åtminstone direkt påverkar varandra.  
Vilken färg har exempelvis b:et i "color yellow color red (a + color green b)", eller vilken storlek har det i "size *4 (a + size / 2 b)"?  
Om man förutsätter en basstorlek på 12, har b:et då storleken 48, 6 eller t o m 24 (vilket skulle kunna gälla som kombination)?  
Numera är detta dock den generella upplösningsregel efter vilken allting ska fungera enhetligt i framtiden.  
Principiellt gäller denna regel för alla grupp-operationer.  
Någon synlig effekt har detta dock bara för teckensnittsattributen, dvs "bold", "ital", "phantom", "size", "color" och "font ":  
Gruppoperationer som har placerats efter varandra behandlas som om var och en av dem skulle vara innesluten av {}.  
De är egentligen kapslade och på varje kapslingssteg finns högst en operation: "size 12 color red font sans size -5 (a + size 8 b)" som "{size 12{color red{font sans{size -5 (a + {size 8 b})}}}} ".  
Sedan tolkas det hela från vänster till höger, varvid en operation genomför de aktuella ändringarna enbart för den tillhörande grupperingen (eller det tillhörande uttrycket).  
De operationer som ligger längre till höger "ersätter" eller "kombineras med "sina föregångare.  
Till dessa hör även deras parenteser samt "super - / subscripts" (upphöjd / nedsänkt skrift), jfr "a + size *2 (b * size -8 c_1)^2 "  
"color..." och "font... "samt "size n" (n är ett decimaltal) ersätter eventuella föregående operationer av samma typ,  
för "size +n", "size -n", "size *n" och "size / n "kombineras operationernas effekter,  
"size *2 size -5 a" skulle vara den dubbla ursprungliga storleken minus 5  
"font sans (a + font serif b)"  
"size *2 (a + size / 2 b)"  
När det gäller StarSymbol-Unicode-Font finns det 2 undantag från dessa regler:  
Detta teckensnitt ignorerar "font "-instruktioner.  
I annat fall skulle man ofta ha andra tecken än de önskade, t ex "font sans (a oplus b)" skulle då varken ha parenteser eller något "oplus ".  
"ital"-instruktionerna ignoreras, t ex "ital (a + b)".  
Detta sker eftersom kursiva matematiska symboler inte är brukliga; inte ens i kombination med kursiv text.  
Dessa kan Du lätt använda i olika sammanhang.  
Du kan använda kommandona Kopiera och Klistra in för att kopiera dem till andra ställen och resultatet är alltid detsamma.  
Dessutom "klarar sig" sådana uttryck bättre när Du ändrar basstorleken på menyn än vad de gör när Du använder "size n ".  
Om Du bara använder "size *" och "size / "(t ex "size *1.24 a eller size / 0.86 a"), bör Du behålla proportionerna.  
Exempel (med basstorlek 12 och 50% för index):  
Fullständigt lika proportioner för "size 18 a_n" och "size *1.5 a_n ".  
I andra sammanhang förhåller det sig dock annorlunda: "x^{size 18 a_n}" och "x^{size *1.5 a_n} "  
Exempel med size +n som jämförelse.  
De ser identiska ut:  
a_{ size 8 n}  
a_{ size +2 n}  
a_{ size *1.333 n}  
Följande exempel ser däremot inte identiska ut:  
x^{ a_{size 8 n}}  
x^{ a_{size +2 n}}  
x^{ a_{size *1.333 n}}  
Tänk på att alla n har olika storlek här.  
Storleken 1.333 fås ur 8 / 6, som är den önskade storleken genom standard-indexstorleken 6. (indexstorlek 50% vid basstorlek 12)  
Index och exponenter  
Här får Du grundläggande information om index och exponenter i %PRODUCTNAME Math.  
De exempel som beskrivs här kan Du utföra själv och på så vis fördjupa Dig mer i detalj. (Citattecknen används bara för att framhäva delar av texten och ingår inte i exemplen.)  
Index och exponent vid ett tecken visas ovanpå varandra, närmare bestämt vänsterjusterat vid bastecknet, t ex a_2^3 "eller ?a^3_2.  
Ordningsföljden har ingen betydelse.  
I stället för '_' och '^ 'kan Du som tidigare använda 'sub' och 'sup '.  
Däremot kan Du inte längre göra på följande sätt:  
a_2_3  
a^2^3  
a_2^3_4  
Varje position för upphöjt / nedsänkt index vid ett bastecken kan bara användas en gång.  
Du måste visa vad Du önskar genom parenteser.  
Följande exempel illustrerar detta:  
a_{ 2_3}  
a^{ 2^3}  
a_2^{ 3_4}  
a_{ 2^3}^{4_5}  
I motsats till andra formelredigerare, där "_" och "^" bara syftar på nästa tecken (alltså vid "a_24 "bara på 2:an), syftar %PRODUCTNAME Math på hela talet / namnet / texten.  
Om Du däremot uttryckligen önskar att den upphöjda och nedsänkta skriften ska stå efter varandra, så skriver Du detta på följande sätt: a_2{ }^3 respektive a^3{ }_2  
Om Du ska skriva tensorer har Du mycket att välja på i %PRODUCTNAME Math.  
Förutom skrivsättet "R_i{}^{jk}{}_l" som även förekommer i andra program, finns det ytterligare alternativ, nämligen "R_i{}^jk{}_l "och "{{R_i}^jk}_l".  
Även upphöjd och nedsänkt index till vänster om bastecknet kan visas, närmare bestämt högerjusterat.  
Till detta används de nya kommandona "lsub" och "lsup ".  
Båda ger exakt samma effekt som "sub" och "sup", men nu till vänster om bastecknet, jfr "a lsub 2 lsup 3 ".  
Reglerna om parentesers entydighet och nödvändighet gäller analogt.  
I princip kan Du även åstadkomma detta med {}_2^3 a.  
Kommandona "sub" och "sup "är även tillgängliga som "rsub" och "rsup ".  
Med dessa alternativ kan Du bl a placera nukleon-, proton - och laddningstal vid kemiska element: "font sans Zn lsub 30 lsup 63 rsup {2+{}}".  
Med kommandona "csub" och "csup "kan Du placera upphöjda och nedsänkta index direkt över respektive under ett tecken, jfr "a csub y csup x".  
Det är även möjligt att ha alla typer av index och exponenter gemensamt: "abc_1^2 lsub 3 lsup 4 csub 55555 csup 66666".  
De flesta enställiga och binära operatorer kan förses med upphöjda och nedsänkta index.  
Här följer två exempel: "a div_2 b a<csub n b +_2 h" och "a toward csub f b x toward csup f y ".  
När Du skriver exempel i kommandofönstret manuellt bör Du tänka på att de befintliga blankstegen är absolut nödvändiga för att exemplet ska byggas upp korrekt.  
Attributegenskaper  
På den här sidan hittar du mer information om attributens egenskaper i %PRODUCTNAME Math. (Citattecknen används bara för att framhäva delar av texten och är inte en del av exemplen eller kommandona.)  
Attributen acute, bar, breve, check, circle, dot, ddot, dddot, grave, hat, tilde och vec har generellt en fast storlek och blir inte bredare (längre) när de står över en lång symbol (jfr t ex dot v och dot vvvvvvv_22222 med det gamla och det nya skrivsättet).  
Som standard centreras de i mitten (jfr dot v_maximum med {dot v}_maximum)  
De enda attribut som fortfarande växer med symbolens längd är "overline", "underline" och "overstrike". ("overstrike "placerar förresten ett streck vågrätt genom "a:et" och inte över a:et.)  
Skillnaderna mellan "bar" och "overline "är viktiga.  
Medan "bar a" och "overline a "fortfarande ser rätt lika ut (förutom att strecket är något kortare hos "bar"), ser de mycket olika ut vid långa symboler.  
Dessa skillnader blir tydliga om Du jämför "bar aaaaa" med "overline aaaaa ".  
Medan strecket hos "bar" bara står över ett tecken, så anpassar sig "overline "till teckenföljdens längd och står således i exemplet över alla fem a.  
Hos vissa teckenuppsättningar kan det t ex förekomma att en linje som infogats med "underline" står för tätt intill bokstaven.  
I ett sådant fall kan Du ta hjälp av en tom grupp, som följande exempel visar.  
Teckensnittet är Times New Roman och bokstaven versalt Q: "underline Q sub {}" i stället för "underline Q ".  
Skalning  
Här finns mer information om skalning i %PRODUCTNAME Math och tillhörande exempel. (Citattecknen används bara för att framhäva delar av texten och ingår inte i exemplen.)  
Fakultetstecknet skalas inte, jfr "fact stack{a#b}" och "fact {a over b} ", utan justeras mot baslinjen eller argumentets mitt.  
Parenteser har generellt också en fast storlek.  
Detta gäller för alla symboler som kan användas som parenteser, jfr "(((a)))"," (stack{a#b#c})", "(a over b) ".  
Parenteser som inleds med "left" respektive "right "anpassas dock alltid till argumentet, jfr "left(left(left(a right)right)right)", "left(stack{a#b#c}right)", "left(a over b right)".  
En del attribut har fasta storlekar och ändrar inte dessa när de står över en lång symbol.  
Du får alltså inte utelämna blankstegen vid inmatning i kommandofönstret.  
Referens  
I den här referensen hittar du alla operatorer, funktioner, symboler och formateringsmöjligheter som är tillgängliga i %PRODUCTNAME Math.  
Många av de kommandon som visas kan du infoga med symbolerna i fönstret Urval eller via snabbmenyn i kommandofönstret.  
Unära och binära operatorer  
Kommandoknapp i urvalsfönstret  
Visning av kommandot i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Unär operator  
Förtecken (+)  
Unär operator  
Förtecken (-)  
Unär operator  
Plusminus (+ -)  
Unär operator  
Minusplus (-+)  
Unär operator  
Logiskt "Inte" (neg)  
Binär operator  
Addition (+)  
Binär operator  
Multiplikation (*)  
Binär operator  
Multiplikation, litet multiplikationstecken (cdot)  
Binär operator  
Multiplikation (times)  
Binär operator  
Subtraktion (-)  
Binär operator  
Division / Bråk (over)  
Binär operator  
Division (div))  
Binär operator  
Division (/)  
Binär operator  
Logisk och-operator (and eller &)  
Binär operator  
Logisk eller-operator (or eller _BAR_)  
Binär operator  
Kedjning av ikoner (circ)  
Binär operator  
Snedstreck / mellan två tecken, varav det vänstra är upphöjt och det högra nedsänkt (wideslash)  
Binär operator  
Snedstreck\ mellan två tecken, varav det högra är upphöjt och det vänstra nedsänkt (widebslash)  
Binär operator  
Additionstecken i cirkel (oplus)  
Binär operator  
Subtraktionstecken i cirkel (ominus)  
Binär operator  
Litet multiplikationstecken i cirkel (odot)  
Binär operator  
Multiplikationstecken times i cirkel (otimes)  
Binär operator  
Snedstreck / i cirkel (odivide)  
Unär operator  
Användardefinierad operator (uoper)  
Binär operator  
Funktionsplatshållare, användardefinierad operator (boper)  
Relationer  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Relation  
Ekvation (=)  
Relation  
Inte lika med (<> eller neq)  
Relation  
Är ungefär (approx)  
Relation  
delar (divides), t.ex. 5 divides 30  
Relation  
delar inte (ndivides), t.ex. 7 ndivides 30  
Relation  
Är mindre än (gt eller <)  
Relation  
Är större än (gt eller >)  
Relation  
Liknar eller är lika med (simeq)  
Relation  
Är parallell med (parallel)  
Relation  
Är ortogonal med (ortho)  
Relation  
Är mindre än eller lika med (leslant)  
Relation  
Är större än eller lika med (geslant)  
Relation  
Liknar (sim)  
Relation  
är identisk / kongruent med (equiv)  
Relation  
Är mindre än eller lika med (le eller <=)  
Relation  
Är större än eller lika med (ge eller >=)  
Relation  
Är proportionell (prop)  
Relation  
strävar mot (toward)  
Operator / logik  
Pil med dubbelstreck åt vänster (dlarrow)  
Operator / logik  
Pil med dubbelstreck åt vänster och höger (dlrarrow)  
Operator / logik  
Pil med dubbelstreck åt höger (drarrow)  
Relation  
Är mycket större än (>> eller gg)  
Relation  
Är mycket mindre än (<< eller ll)  
Binär operator / Relation  
är definierad som / definitionsmässigt lika med (def)  
Relation  
Korrespondenstecken bild från (transl)  
Relation  
Korrespondenstecken original från (transr)  
Mängdoperatorer  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Mängdoperator  
tillhör (in)  
Mängdoperator  
tillhör inte (notin)  
Mängdoperator  
Innehåller (owns eller ni)  
Matematisk symbol  
Tomma mängden (emptyset)  
Mängdoperator  
Genomsnitt av mängder (intersection)  
Mängdoperator  
Union av mängder (union)  
Mängdoperator  
Differensmängd (setminus eller bslash)  
Mängdoperator  
Snedstreck / för kvot (slash) mellan tecken, t ex A slash B slash C  
Matematisk symbol  
Kardinaltal (aleph)  
Mängdoperator  
Delmängd (subset)  
Mängdoperator  
Delmängd eller lika med (subseteq)  
Mängdoperator  
Grundmängd (supset)  
Mängdoperator  
Grundmängd eller lika med (supseteq)  
Mängdoperator  
ej delmängd av (nsubset)  
Mängdoperator  
Ej delmängd eller lika med (nsubseteq)  
Mängdoperator  
ej grundmängd (nsupset)  
Mängdoperator  
Ej grundmängd eller lika med (nsupseteq)  
Matematisk symbol  
naturligt tal (setn)  
Matematisk symbol  
heltal (setz)  
Matematisk symbol  
rationellt tal (setq)  
Matematisk symbol  
reellt tal (setr)  
Matematisk symbol  
komplext tal (setc)  
Funktioner  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Funktion  
Naturlig exponentialfunktion (func e^{})  
Funktion  
Naturlig logaritm (ln)  
Funktion  
Allmän exponentialfunktion (exp)  
Funktion  
Allmän logaritm (log)  
Funktion / binär operator  
n:te potensen av x (sup)  
Funktion  
Sinus (sin)  
Funktion  
Cosinus (cos)  
Funktion  
Tangens (tan)  
Funktion  
Cotangens (cot)  
Funktion  
Kvadratrot (sqrt)  
Funktion  
Arcussinus (arcsin)  
Funktion  
Arcuscosinus (arccos)  
Funktion  
Arcustangens (arctan)  
Funktion  
Arcuscotangens (arccot)  
Funktion  
n:te kvadratroten ur x( nroot)  
Funktion  
Sinus hyperbolicus (sinh)  
Funktion  
Cosinus hyperbolicus (cosh)  
Funktion  
Tangens hyperbolicus (tanh)  
Funktion  
Cotangens hyperbolicus (coth)  
Funktion  
Absolutvärde (abs)  
Funktion  
Area sinus hyperbolicus (arsinh)  
Funktion  
Area cosinus hyperbolicus (arcosh)  
Funktion  
Area tangens hyperbolicus (artanh)  
Funktion  
Area cotangens hyperbolicus (arcoth)  
Funktion  
Fakultet (fact)  
Matematisk symbol  
Omvänt epsilon (backepsilon)  
Binär operator  
x med index n (sub)  
Operatorer  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Operator  
Limes (lim)  
Operator  
Summa (sum)  
Operator  
Produkt (prod)  
Operator  
Koprodukt (coprod)  
Operator  
Områdesuppgift från... till (from to)  
Operator  
Integral (int)  
Operator  
Dubbelintegral (iint)  
Operator  
Tredubbel integral (iiint)  
Operator  
En operators nedre gräns (from)  
Operator  
Kurvintegral (lint)  
Operator  
dubbel kurvintegral (llint)  
Operator  
tredubbel kurvintegral (lllint)  
Operator  
En operators övre gräns (to)  
Operator  
Limes inferior (liminf)  
Operator  
Limes superior (limsup)  
Operator  
Platshållare, användardefinierad operator (oper)  
Attribut  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Attribut med fast teckenbredd  
Accent åt höger ovanför ett tecken (acute)  
Attribut med fast teckenbredd  
Accent åt vänster (grave) ovanför ett tecken  
Attribut med fast teckenbredd  
omvänt tak (check)  
Attribut med fast teckenbredd  
"Omvänt tak" ovanför ett tecken (breve)  
Attribut med fast teckenbredd  
Cirkel ovanför ett tecken (circle)  
Attribut med fast teckenbredd  
Vektorpil ovanför ett tecken (vec)  
Attribut med fast teckenbredd  
Tilde ovanför ett tecken (tilde)  
Attribut med fast teckenbredd  
"Tak" ovanför ett tecken (hat)  
Attribut med fast teckenbredd  
Vågrätt streck över ett tecken (bar)  
Attribut med fast teckenbredd  
Punkt ovanför ett tecken (dot)  
Attribut med variabel teckenbredd  
bred vektorpil som anpassar sig till teckenstorleken (widevec)  
Attribut med variabel teckenbredd  
brett tilde, som anpassar sig till teckenstorleken (widetilde)  
Attribut med variabel teckenbredd  
brett tak, som anpassar sig till teckenstorleken (widehat)  
Attribut med fast teckenbredd  
Två punkter ovanför ett tecken (ddot)  
Attribut med variabel teckenbredd  
Vågrätt streck över ett tecken (overline)  
Attribut med variabel teckenbredd  
Vågrätt streck under ett tecken (underline)  
Attribut med variabel teckenbredd  
Vågrätt streck genom ett tecken (overstrike)  
Attribut med fast teckenbredd  
Tre punkter ovanför ett tecken (dddot)  
Teckenattribut  
Fantomtecken (phantom)  
Teckenattribut  
Fet (bold)  
Teckenattribut  
Kursiv (ital)  
Teckenattribut, ändra storlek  
Storleksangivelserna kan förses med argument i form av n, +n, -n *n eller / n.  
En procentuell förändring med t ex 17% anges i formen *1,17.  
Teckenattribut, ändra teckensnitt  
Först anger du teckensnittets namn, sans, serif eller fixed, och därefter de tecken som ska ändras.  
Teckenattribut  
Först anger du färgens namn (black, white, cyan, magenta, red, blue, green och yellow), och därefter de tecken som ska ändras.  
Färgattribut måste anges direkt i kommandofönstret.  
Teckenattribut  
Upphäva attributet kursiv (nitalic)  
Teckenattribut  
Upphäva attributet fet (nbold)  
Övrigt  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Matematisk symbol  
Oändlig (infinity eller infty)  
Matematisk symbol  
Partiell derivata eller också en mängds begränsning (partial)  
Matematisk symbol  
Nablavektor (nabla)  
Operator / logik  
Existenskvantifikator, det finns minst en (exists)  
Operator / logik  
Allkvantifikator, för alla (forall)  
Operator / fysik  
h med vågrätt streck (hbar)  
Operator / fysik  
Lambda med vågrätt streck (lambdabar)  
Matematisk symbol  
Realdelen av ett komplext tal (re)  
Matematisk symbol  
Imaginärdelen av ett komplext tal (im)  
Matematisk symbol  
p-funktion (wp), Weierstrass p  
Operator  
Pil till vänster (leftarrow)  
Operator  
Pil till höger (rightarrow)  
Operator  
Pil uppåt (uparrow)  
Operator  
Pil nedåt (downarrow)  
Annan symbol  
Tre prickar vågrätt nere (dotslow)  
Annan symbol  
Tre prickar vågrätt i teckenmitten (dotsaxis)  
Annan symbol  
Tre prickar diagonalt nerifrån vänster och upp till höger (dotsup eller dotsdiag)  
Annan symbol  
Tre prickar lodrätt (dotsvert)  
Annan symbol  
Tre prickar diagonalt uppifrån vänster och ned till höger (dotsdown)  
Annan symbol  
Platshållare <?>  
Parenteser  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Parentes med grupperingsfunktion  
Normal rund vänster och höger parentes  
Parentes med grupperingsfunktion  
Vänster och höger hakparentes  
Parentes med grupperingsfunktion  
Dubbel vänster och höger hakparentes (ldbracket... rdbracket)  
Parentes med grupperingsfunktion  
Vänster och höger lodrät linje (lline... rline)  
Parentes med grupperingsfunktion  
Dubbel vågrät vänster - och högerlinje (ldline... rdline)  
Parentes med grupperingsfunktion  
Vänster och höger klammerparentes, mängdparentes (lbrace... rbrace)  
Parentes med grupperingsfunktion  
Vänster och höger vinkelparentes (langle... rangle)  
Parentes med grupperingsfunktion  
Vänster och höger vinkelparentes för operator (langle... mline...rangle)  
Parentes med grupperingsfunktion  
Vänster och höger grupparentes.  
De visas inte i dokumentet och behöver ingen plats.  
se normala parenteser  
Parentes med grupperingsfunktion  
Automatisk storleksanpassning i parenteserna genom placering av left och right framför (left... right...), t ex left(a over b right) eller left lceil... right lceil.  
På detta sätt kan Du ändra runda parenteser, hakparenteser, dubbla hakparenteser, enkla parenteser, dubbla enkla parenteser, klammerparenteser, vinkelparenteser och operator-parenteser.  
se hakparenteser  
Parentes med grupperingsfunktion, skalbar  
Skalbara hakparenteser, i kommandofönstret sker inmatningen enligt mönstret (left[... right]).  
se dubbla hakparenteser  
Parentes med grupperingsfunktion, skalbar  
Dubbla skalbara hakparenteser, (left ldbracket... right rdbracket)  
se lodräta parenteser  
Parentes med grupperingsfunktion, skalbar  
Mängdparenteser, (mata in left lbrace... right rbrace)  
se dubbla lodräta parenteser  
Parentes med grupperingsfunktion, skalbar  
Enkla skalbara linjer, (left lline... right rline)  
se klammerparenteser  
Parentes med grupperingsfunktion, skalbar  
Dubbla skalbara linjer, (left ldline... right rdline)  
se vinkelparenteser  
Parentes med grupperingsfunktion, skalbar  
Skalbara vinkelparenteser, (left langle... right rangle)  
se operatorparenteser  
Parentes med grupperingsfunktion  
Skalbar vänster och höger vinkelparentes för operator (left langle... mline...right rangle)  
Parentes med grupperingsfunktion  
Skalbara klammerparenteser uppe (... overbrace...)  
Parentes med grupperingsfunktion  
Skalbara klammerparenteser nere (... underbrace...)  
Parentes med grupperingsfunktion  
Vänster och höger linje med kanter nere (lfloor... rfloor)  
Parentes med grupperingsfunktion  
Vänster och höger linje med kanter uppe (lceil... rceil)  
se klammerparenteser  
Parentes, också fristående, utan grupperingsfunktion  
Vänster klammerparentes: \lbrace eller \{ resp. rcchte klammerparentes: \rbrace eller\})  
se normala parenteser  
Parentes, också fristående, utan grupperingsfunktion  
Vänster och höger parentes: \( eller\)  
se hakparenteser  
Parentes, också fristående, utan grupperingsfunktion  
Vänster och höger hakparentes: \[ eller\]  
se vinkelparenteser  
Parentes, också fristående, utan grupperingsfunktion  
Vänster och höger vinkelparentes: \langle eller \rangle  
se lodrät linje  
Parentes, också fristående, utan grupperingsfunktion  
Vänster och höger lodrät linje: \lline eller \rline  
se dubbel lodrät linje  
Parentes, också fristående, utan grupperingsfunktion  
Dubbel vänster och höger linje: \ldline eller \rdline  
se linje med kanter nere  
Parentes, också fristående, utan grupperingsfunktion  
Vänster och höger linje med kanter nere: \lfloor eller \rfloor  
se linje med kanter uppe  
Parentes, också fristående, utan grupperingsfunktion  
Vänster och höger linje med kanter uppe: \lceil eller \rceil  
Formateringar  
Kommandoknapp i urvalsfönstret  
Visning av kommando i en formel  
Grupp  
Betydelse (inom parentes: kommando i kommandofönstret)  
Index o. exponenter (sub - och superscript)  
Vänster exponent (lsup)  
Index o. exponenter (sub - och superscript)  
Exponent direkt ovanför ett tecken (csup)  
Index o. exponenter (sub - och superscript)  
Höger exponent (^ eller sup eller rsup)  
Formatering  
Binom (binom)  
Formatering  
Ny rad (newline)  
Index o. exponenter (sub - och superscript)  
Vänster index (lsub)  
Index o. exponenter (sub - och superscript)  
Index direkt under ett tecken (csub)  
Index o. exponenter (sub - och superscript)  
Höger index (_ eller sub eller rsub)  
Formatering  
Stack (stack) anges enligt mönstret: stack{x#y#z}  
Formatering  
Litet mellanrum / Litet blanksteg (')  
Formatering  
Horisontell justering (alignl eller alignc eller alignr)  
Formatering  
Horisontell justering centrerat (alignc)  
Formatering  
Horisontell justering till höger (alignr)  
Formatering  
Matris (matrix), anges enligt mönstret: matrix{a#b##c#d}  
Formatering  
Stort mellanrum / blanksteg (~)  
Övrigt  
Välj bland diverse matematiska symboler när du ska bygga upp en %PRODUCTNAME Math -formel.  
Du hittar alla tillgängliga operatorer om du öppnar snabbmenyn i fönstret Kommandon och sedan välja Övrigt.  
Symboler som inte kan skapas via urvalsfönstret eller snabbmenyn måste du skriva in direkt i kommandofönstret.  
Du kan naturligtvis också bygga upp alla andra symboler manuellt.  
Symbolerna i detalj:  
Med ikonen infogar du en partiell differential eller en mängds begränsning.  
Du kan också skriva partial direkt i kommandofönstret.  
Partial  
Med ikonen infogar du tecknet för oändlig.  
Du kan även skapa tecknet genom att skriva infinity eller infty i kommandofönstret.  
Oändlig:  
Med ikonen infogar du Nablavektorn.  
I stället för att använda ikonen kan du skriva nabla direkt i kommandofönstret.  
Nabla  
Med ikonen infogar du existenskvantifikatorn "det finns".  
I stället för att använda ikonen kan du skriva exists direkt i kommandofönstret.  
Det finns  
Med ikonen infogar du allkvantifikatorn "för alla".  
I stället för att använda ikonen kan du skriva forall direkt i kommandofönstret.  
För alla  
Med ikonen infogar du den lilla bokstaven h med ett vågrät streck.  
I stället för att använda ikonen kan du skriva hbar direkt i kommandofönstret.  
Strukna h  
Med ikonen infogar du den lilla grekiska bokstaven lambda med ett vågrät streck.  
I stället för att använda ikonen kan du skriva lambdabar direkt i kommandofönstret.  
Strukna lambda  
Med ikonen infogar du tecknet för ett komplext tals realdel.  
Du kan också ange kommandot re, vilket ger samma resultat.  
Realdel  
Med ikonen infogar du tecknet för ett komplext tals imaginärdel.  
I stället för att använda ikonen kan du ange kommandot im direkt.  
Imaginärdel  
Med ikonen infogar du ett Weierstrass p.  
Du kan också infoga p-funktionen direkt genom att ange wp i kommandofönstret.  
Weierstrass p  
Med ikonen infogar du en vänsterpil.  
Du uppnår samma resultat genom att skriva leftarrow.  
Pil åt vänster  
Med ikonen infogar du en högerpil.  
Du kan också skapa en sådan genom att skriva rightarrow i kommandofönstret.  
Pil åt höger  
Med ikonen infogar du en uppåtpil.  
Du kan också skriva uparrow direkt i kommandofönstret.  
Pil uppåt  
Med ikonen infogar du en nedåtpil.  
Du uppnår samma resultat genom att skriva downarrow.  
Pil nedåt  
Med ikonen infogar du tre vågräta punkter nedtill.  
I stället för att använda ikonen kan du också skriva dotslow direkt i kommandofönstret.  
Punkter nere  
Med ikonen infogar du tre vågräta punkter i höjd med teckenmitten.  
I stället för att använda ikonen kan du ange kommandot dotaxis direkt i kommandofönstret.  
Punkter i mitten  
Med ikonen infogar du tre lodräta punkter.  
I stället för att använda ikonen kan du också skriva dotsvert direkt i kommandofönstret.  
Punkter vertikalt  
Med ikonen infogar du tre punkter på diagonalen nerifrån vänster upp till höger.  
I stället för att använda ikonen kan du också skriva dotsup eller dotsdiag direkt i kommandofönstret.  
Punkter uppåt  
Med ikonen infogar du tre punkter som löper diagonalt uppifrån vänster och ner till höger.  
I stället för att använda ikonen kan du också skriva kommandot dotsdown direkt i kommandofönstret.  
Punkter nedåt  
Du infogar ett omvänt epsilon genom att mata in backepsilon i kommandofönstret.  
Det här kommandot är inte tillgängligt via Övrigt -menyn.  
Om du vill infoga en platshållare i ditt dokument matar du in <?> i kommandofönstret.  
Kommandot är inte tillgängligt via Övrigt -menyn.  
Teckensnitt  
Här definierar du de teckensnitt som används för vissa formelelement.  
Formelteckensnitt  
I det här området definierar Du teckensnitten för de formelelement som Du infogar med %PRODUCTNAME, dvs för variabler, funktioner och tal.  
Här väljer Du även teckensnitt för de texter som Du infogar.  
I listrutorna visas först bara de förinställda teckensnitten för varje område.  
Efter posten Funktioner kan Du t ex bara välja teckensnittet Times New Roman.  
Om Du alltid, eller emellanåt, vill visa funktionerna med ett annat teckensnitt, kan Du utöka listrutan med ytterligare teckensnitt, som Du sedan kan välja bland.  
Om Du vill utöka urvalet i listrutan, använder Du kommandoknappen Ändra.  
Om Du vill framhäva enstaka textdelar med något annat teckensnitt än det som definierats för alla texter, så definierar Du detta med kommandot FONT i kommandofönstret.  
Variabler  
Här väljer Du teckensnitt för variablerna i formeln.  
I formeln x=SIN( y) är x och y variabler.  
Funktioner  
Här väljer Du teckensnitt för funktionernas namn och övriga delar.  
I formeln x=SIN( y) är detta tecknen =SIN ().  
Tal  
Här väljer Du teckensnitt för talen i formeln.  
Text  
Här väljer Du teckensnitt för alla övriga texter i formeln.  
Användarteckensnitt  
I det här området definierar Du tre teckensnitt med vilka Du kan formatera andra textdelar i formeln.  
Tillgängliga alternativ är de tre basteckensnitten Serif, Sans och Fixed.  
Till varje basteckensnitt som installerats som standard kan Du lägga till ytterligare ett valfritt.  
Du kan välja vilket teckensnitt som helst, förutsatt att det har installerats i systemet.  
Om Du vill utöka urvalet i listrutorna, använder Du kommandoknappen Ändra.  
Dessa användarteckensnitt används om Du anger ett annat teckensnitt i kommandofönstret med kommandot FONT.  
Du kan testa detta genom att kopiera följande text till kommandofönstret:  
font sans "Vi presenterar:" newline  
font serif "%PRODUCTNAME Math," newline  
font serif "formel-editorn i" newline  
font sans "%PRODUCTNAME %PRODUCTVERSION" newline  
font serif "som levereras av" newline  
font fixed "Sun Microsystems"  
Serif  
Här väljer Du det teckensnitt som ska användas för formateringen font serif i formeln.  
Seriffer är de små "tvärstreck" som t ex visas nedtill på ett versalt A i ett seriffteckensnitt som Times.  
De förbättrar läsbarheten i löpande text.  
Sans  
Här väljer Du det teckensnitt som ska användas för formateringen font sans i formeln.  
Teckensnitt utan seriffer (sans serif), som t ex Arial, används ofta för överskrifter.  
Fixed  
Här väljer Du det teckensnitt som ska användas för formateringen font fixed i formeln.  
Icke-proportionella teckensnitt som Courier kan Du med fördel använda i tabeller.  
Ändra  
Klicka på den här knappen om Du vill öppna dialogrutan Teckensnitt, där Du kan definiera teckensnitt och attribut för de enskilda formel - och användarteckensnitten.  
När Du klickar på den här kommandoknappen visas först en popupmeny i vilken Du kan välja område.  
Standard  
Om Du klickar på den här kommandoknappen, sparas de gjorda ändringarna som standard för alla nya formler.  
Innan ändringarna sparas får Du en kontrollfråga.  
Teckensnitt  
I den här dialogrutan väljer Du ett teckensnitt som sedan är tillgängligt för det valda området i dialogrutan Teckensnitt.  
Teckensnitt  
I det här kombinationsfältet anger Du önskat teckensnitt.  
Ange det exakta namnet.  
Du kan också välja bland de teckensnitt som är tillgängliga i systemet i listrutan nedanför.  
Klicka på det önskade teckensnittet.  
Exempel  
Här presenteras en förhandsvisning av det valda teckensnittet med dess attribut.  
Attribut  
I det här området kan Du tilldela det valda teckensnittet ytterligare attribut.  
Fet  
Om Du markerar den här kryssrutan visas teckensnittet fetstilt.  
Kursiv  
Om Du markerar den här kryssrutan visas teckensnittet kursivt.  
Teckenstorlekar  
I den här dialogrutan definierar du teckenstorlekarna i formeln.  
Du väljer en basstorlek och definierar alla element i formeln i procentuell relation till basen.  
Basstorlek  
Här väljer du den basstorlek till vilken alla andra storlekar relaterar.  
I det här rotationsfält et kan du använda enheten punkt (pt, point) eller någon annan enhet som programmet sedan räknar om till pt.  
Om du vill ändra den använda standardstorleken (12 pt) som används i %PRODUCTNAME Math, så måste du först ställa in den nya storleken (t.ex. 11 pt) i rotationsfältet Basstorlek och sedan klicka på kommandoknappen Standard.  
Relativa storlekar  
I det här området väljer Du de relativa storlekarna i förhållande till basstorleken.  
Text  
Här väljer Du textens relativa storlek.  
Som standard är den 100%.  
Index  
Här väljer Du relativ storlek för index.  
Som standard är den 50%.  
Funktioner  
Här väljer Du relativ storlek för funktionernas namn och övriga element.  
Som standard är den 100%.  
Operatorer  
Här väljer Du relativ storlek för de matematiska operatorerna.  
Som standard är den 100%.  
Gränser  
Här väljer Du relativ storlek för gränserna, t ex under och över summatecknen.  
Som standard är den 50%.  
Standard  
Om Du klickar på den här kommandoknappen, sparas de gjorda ändringarna som standard för alla nya formler.  
Innan ändringarna sparas får Du en kontrollfråga.  
Avstånd  
I den här dialogrutan definierar du avstånd för formelelement, t.ex. index, gränser, operatorer.  
Du anger avstånden i procent, i relation till den basstorlek som du har valt i Format - Teckenstorlekar.  
Även värden på 0% och över 100% är möjliga.  
Med kommandoknappen Kategori väljer Du de formelelement för vilka Du ska definiera avstånd.  
Dialogrutan ändras så att dess utseende motsvarar den valda kategorin.  
I ett förhandsvisningsfönster visas vilka avstånd Du kan ändra i de aktuella rotationsfälten.  
Du kan välja bland följande kategorier:  
Avstånd, Index, Bråk, Bråkstreck, Gränser, Parenteser, Matriser, Ornament, Operatorer och Marginaler.  
Kategori  
När Du har klickat på den här kommandoknappen, kan Du välja den kategori vars avstånd Du vill bestämma.  
Avstånd  
Här bestämmer Du avstånden mellan variabler och operatorer, mellan rader och mellan rottecken och det tal varur roten ska dras.  
Avstånd  
Här definierar Du avståndet mellan variabler och operatorer.  
Radavstånd  
Här definierar Du avståndet mellan rader.  
Rotavstånd  
Här definierar Du avståndet mellan rottecken och det tal varur roten ska dras.  
Index  
Här definierar Du avståndet för upphöjda och nedsänkta index.  
Upphöjning  
Här definierar Du avståndet för upphöjda index.  
Nedsänkning  
Här definierar Du avståndet för nedsänkta index.  
Bråk  
Här definierar Du avståndet mellan bråkstreck och täljare eller nämnare.  
Täljare, höjd  
Här definierar Du avståndet mellan bråkstreck och täljare.  
Nämnare, djup  
Här definierar Du avståndet mellan bråkstreck och nämnare.  
Bråkstreck  
Här definierar Du bråkstreckens överskjutning och linjestyrka.  
Överskjutning  
Här definierar Du bråkstreckens överskjutning.  
Linjestyrka  
Här definierar Du bråkstreckens linjestyrka.  
Gränser  
Här definierar Du avstånden mellan t ex summatecken och gränsvillkor.  
Gränshöjd  
Här definierar Du avståndet mellan summatecken och övre gräns.  
Gränsdjup  
Här definierar Du avståndet mellan summatecken och startvillkor.  
Parenteser  
Här definierar Du avstånden mellan stora parenteser och deras innehåll.  
Vänster / höger överstorlek  
Här definierar Du det vertikala avståndet mellan parentesinnehållets överkant och parentesens övre slut.  
Avstånd  
Här definierar Du det horisontella avståndet mellan parentesinnehållet och parentesens övre slut.  
Skala alla parenteser  
Om du markerar den här rutan, så skalas alla parentestyper.  
Om du sedan skriver t.ex. (a over b) i kommandofönstret, så omfattar parenteserna argumentets hela höjd.  
En sådan effekt uppnår du normalt bara om du skriver left (a over b right).  
Överstorlek  
I det här rotationsfältet anger du den procentuella överstorlek som parenteserna ska ha i förhållande till sitt innehåll.  
Vid 0 procent är parenteserna satta så att de omsluter argumentet ungefär i samma höjd.  
Ju högre det inställda värdet är, desto större blir det lodräta avståndet mellan parentesinnehållet och parentesernas utvändiga marginal.  
Du kan bara använda rutan i kombination med Skala alla parenteser.  
Genom att kombinera dessa inställningar kan du lätt bygga upp växande kapslade parenteser.  
Ange t.ex. 5 procent för Vänster / höger överstorlek.  
Markera rutan Skala alla parenteser och ange 0 procent i det tillhörande rotationsfältet Överstorlek.  
Resultatet ser du om du skriver följande kapslingar: left (left (left ((((a over b))) right) right) right)  
Matriser  
Här definierar Du de avstånd som element i matriser har till varandra.  
Radavstånd  
Här definierar Du matriselementens radavstånd.  
Kolumnavstånd  
Här definierar Du matriselementens kolumnavstånd.  
Ornament  
Här definierar Du de avstånd som ornamenten har till variablerna.  
Primärhöjd  
Här definierar Du ornamentens höjd över baslinjen.  
Minimiavstånd  
Här definierar Du ornamentens minimiavstånd över variablerna.  
Om Du vill placera flera vågräta streck över ett tecken, t ex overline {overline A intersection overline B}, och om avståndet mellan strecken är för litet, kan Du öka detta i rotationsfältet Minimiavstånd.  
Ange helt enkelt ett högre procentvärde.  
Operatorer  
Här definierar Du avstånden mellan operatorer och variabler eller tal.  
Överstorlek  
Här definierar Du den extra höjd som operatorernas överkant har över variablerna.  
Avstånd  
Här definierar Du det horisontella avståndet mellan operatorer och variabler.  
Marginaler  
Här kan Du göra marginalinställningar för formeln.  
Detta alternativ är särskilt intressant om Du t ex ska infoga formeln i texter i %PRODUCTNAME Writer.  
Se till att Du inte anger 0 som storlek.  
I så fall uppstår naturligtvis problem med visningen i de områden som gränsar till den omgivande texten.  
Vänster  
Här anger Du den vänstra marginalen mellan formel och omgivning.  
Höger  
Här anger Du den högra marginalen mellan formel och omgivning.  
Uppe  
Här anger Du den övre marginalen mellan formel och omgivning.  
Nere  
Här anger Du den undre marginalen mellan formel och omgivning.  
Standard  
Om Du klickar på den här kommandoknappen, sparas de gjorda ändringarna som standard för alla nya formler.  
Innan ändringarna sparas får Du en kontrollfråga.  
Den här "Standard "-kommandoknappens funktion skiljer sig från övriga kommandoknappar med samma namn i %PRODUCTNAME!  
Justering  
Här definierar du justeringen för flerradiga formler och sådana med flera delar på en rad.  
Flerradiga formler får du om du anger kommandot NEWLINE på kommandoraden.  
Men även täljare och nämnare i ett bråk räknas som flerradiga i denna bemärkelse.  
Ett likhetstecken i en formel delar formeln i en vänster - och högerdel (om likhetstecknet inte står i t.ex. ett parentesuttryck).  
Horisontell  
Det här området används för vågrät justering av flerradiga formler.  
Vänster  
Formelraderna placeras vänsterjusterat under varandra.  
Om Du snabbt vill vänsterjustera en viss formelrad, t ex om Du vill tilldela den till en text, så placerar Du helt enkelt två citattecken "" i dess början.  
Den tomma sträng som Du därigenom skapar indikerar för %PRODUCTNAME Math att det är frågan om en textrad.  
Eftersom texter alltid vänsterjusteras, hamnar även formelraden där.  
Alla övriga formler centreras på nytt.  
Om Du däremot vill centrera en text, inleder Du texten med en tom grupp {}.  
Detaljerna anger Du i menyn Format - Avstånd....  
Centrerad  
Formelraderna placeras centrerat under varandra.  
Höger  
Formelraderna placeras högerjusterat under varandra.  
Standard  
Om Du klickar på den här kommandoknappen, sparas de gjorda ändringarna som standard för alla nya formler.  
Innan ändringarna sparas får Du en kontrollfråga.  
Textläge  
Med det här kommandot sätter du på resp. stänger av textläget.  
I textläget visas en formel med samma höjd som en textrad.  
Katalog  
Med det här kommandot öppnar du dialogrutan Symboler.  
I den här dialogrutan väljer du en symbol som ska infogas i formeln.  
Välj ett tecken i dialogrutan och klicka på Överta, så infogas det kommando som visar det här tecknet i kommandofönstret.  
För lilla grekiska alfa är kommandot "%alpha" (bara små bokstäver), och för stora alfa är det "%ALPHA "(enbart versaler).  
Symbolset  
I den här listrutan väljer du ett symbolset som visas i fältet som finns nedanför.  
Symbol  
I det här området visas symbolen och namnet på symbolen.  
Nä du skriver namnet på en symbol i kommandofönstret måste du skriva exakt på det sättet som det är skrivet här när det gäller stora och små bokstäver.  
Redigera...  
Med den här kommandoknappen kommer du till dialogrutan Redigera symboler.  
Redigera symboler  
I den här dialogrutan tilldelar du symbolteckenuppsättningen i %PRODUCTNAME tecken, ändrar symbolbeteckningar eller redigerar hela symbolset.  
Du kan definiera nya symbolset, ge symboler namn och lägga till dem i symbolseten.  
Du kan redigera befintliga symbolset.  
Gammal symbol  
I det här fältet väljer du den aktuella symbolen med dess namn.  
Symbolen visas i det vänstra förhandsvisningsfönstret i dialogrutans nedre del.  
Där visas dessutom namnen på symbolen och symbolsetet.  
Gammalt symbolset  
Här ser du namnet på det aktuella symbolsetet och kan välja ett annat set.  
Symbol  
Här anger du namnet för en ny symbol som ska läggas till, eller ändrar namnet på en symbol.  
Lägga till ny symbol  
Om du vill lägga till ett nytt tecken till ett symbolset, väljer du först ett Teckensnitt och klickar på det önskade tecknet i listrutan.  
Ge symbolen ett namn i fältet Symbol.  
Välj ett symbolset eller ange namnet på ett nytt symbolset.  
Den symbol som ska infogas visas i det högra av de båda förhandsvisningsfönstren.  
Klicka på OK.  
Ändra namn på en symbol  
Skriv sedan det nya namnet i fältet Symbol.  
Kontrollera om det önskade tecknet verkligen visas i förhandsvisningsfönstret innan du klickar på kommandoknappen Ändra.  
Klicka på OK.  
Symbolset  
Du väljer ett set som ska ändras i listan, eller skapar ett nytt genom att ange dess namn.  
Skapa nytt symbolset  
Om du vill skapa ett nytt symbolset anger du ett namn för det i kombinationsfältet Symbolset och lägger till minst en symbol.  
Du stänger dialogrutan med OK.  
Det nya symbolsetet är nu tillgängligt med det nya namnet.  
Teckensnitt  
Ett %PRODUCTNAME Math-symbolset kan innehålla tecken från olika teckensnitt.  
Område  
Om du har valt ett icke-symbol-teckensnitt i fältet Teckensnitt kan du välja ett Unicode-område här.  
Teckenstil  
Välj en annan teckenstil.  
Lägg till  
Om du klickar på den här kommandoknappen så läggs det tecken till som visas i det högra förhandsvisningsfönstret under namnet i fältet Symbol till symbolsetet vars namn står i fältet Symbolset.  
Den här kommandoknappen kan du bara använda om du har skrivit ett nytt namn i fältet Symbol eller i fältet Symbolset.  
Namn får inte tilldelas dubbelt.  
Ändra  
Om du klickar på den här kommandoknappen får symbolen som visas i det vänstra förhandsvisningsfönstret och vars gamla namn står i fältet Gammal symbol ett nytt namn som du har skrivit in i fältet Symbol.  
Flytta symbol till annat symbolset  
Anta att du vill flytta stort ALFA från symbolsetet "Grekiskt" till setet "Special ".  
Välj det gamla setet (Grekiskt) och sedan symbolen ALFA från de båda övre listrutorna.  
Det visas i det vänstra förhandsvisningsfönstret.  
Välj symbolsetet "Special" i kombinationsfältet Symbolset Klicka på Ändra och sedan på OK.  
Symbolen ALFA finns nu bara i symbolsetet "Special"  
Radera  
Med det här kommandot raderar du den symbol som står i det vänstra förhandsvisningsfönstret från det aktuella symbolsetet.  
Du får ingen kontrollfråga.  
Med den sista symbolen i ett symbolset raderar du också symbolsetet.  
Om Du har gjort något misstag kan Du stänga dialogrutan med Avbryt, varvid de gjorda ändringarna inte sparas.  
Importera formel  
Med det här kommandot öppnar du en dialogruta där du kan importera en formel.  
Dialogrutan Infoga är uppbyggd på samma sätt som dialogrutan Öppna på menyn Arkiv.  
Här kan du ladda och redigera en formel som är sparad som fil i kommandofönstret och (när du har valt kommandot Visa - Uppdatera eventuellt) visa den.  
Formelmarkör  
Här sätter du på och stänger av formelmarkören.  
Den del av formeln där inmatningsmarkören står i kommandofönstret markeras med en tunn ram när formelmarkören är aktiverad.  
Du kan också klicka på en del av formeln i dokumentet för att flytta markören i kommandofönstret till motsvarande plats.  
Om du dubbelklickar i dokumentet flyttas markören i kommandofönstret och samtidigt markeras motsvarande ställe.  
Här följer några exempel som visar hur det fungerar:  
Sin (x)  
Alla komponenter markeras av formelmarkören.  
Size *2 bold italic w  
Bara bokstaven w markeras, eftersom de andra tecknen inte visas i textfönstret.  
Sum from a to b x_i^2  
Komponenterna from och to är tecken som inte visas och alltså inte heller markeras.  
"Detta är en text."  
Hela texten inom citattecken markeras.  
<?>  
Alla komponenterna i platshållaren markeras.  
Kortkommandon för formeldokument  
Här hittar du tangentkombinationer som kan förenkla arbetet med formeldokument.  
Dessutom gäller de allmänna tangentkombinationerna i %PRODUCTNAME.  
De kommandon vars tangentkombinationer listas här finns i menyerna Redigera och Visa.  
Tangentkombinationer för funktioner i formeldokument  
Tangentkombination  
Effekt  
F2  
Hoppar till nästa platshållare i kommandofönstret  
Skift+F2  
Hoppar till föregående platshållare  
F3  
Hoppar till nästa fel  
Skift+F3  
Hoppar till föregående fel  
F9  
Uppdaterar visningen  
Justera formeldelar manuellt  
Hur kan tecken i %PRODUCTNAME Math snabbt och lätt justeras?  
Utnyttja möjligheten att definiera tomma grupper och teckensträngar.  
De behöver ingen plats, men innehåller information som hjälper dig vid justeringen.  
Om du vill skapa tomma grupper matar du in klammerparanteser {} i kommandofönstret.  
I följande exempel visas hur man gör en radbrytning där plustecknen står under varandra, trots att ett tecken mindre matas in i den övre raden: a+a+a+{} newline {}{}{}{}{ }a+a+a+a  
De definieras med dubbla citationstecken "".  
Undvik att använda typografiska citationstecken.  
Exempel: "Ett ytterligare exempel." newline a+b newline ""c-d  
Ändra standardattribut  
Går det att ändra standardformateringar i %PRODUCTNAME Math?  
Om delar av en formel i StarMath enligt standard är fett eller kursivt formaterade kan du ändra attributen med kommandona "nbold" och "nitalic ".  
Följande exempel förtydligar detta: nitalic a + bold b.  
I den här formeln visas a inte längre kursivt, b:et får tvärt emot förinställningen attributet fet.  
Plustecknet kan för övrigt inte ändras på det här sättet.  
Sammanfatta formeldelar i parenteser  
Så här matar du in bråk i en formel.  
De sammanhörande värdena måste sammanfattas med en parentes för ett bråk vars täljare eller nämnare består av en produkt, en summa osv.  
Använd följande syntax: "{a + c} over 2 = m" eller "m = {a + c} over 2 "  
Mata in kommentar  
Hur kan en formel förses med kommentarer som inte visas i dokumentet?  
En kommentar börjar med dubbla procenttecken%% och fortsätter till nästa radslutstecken (returtangenten).  
Allt som står däremellan ignoreras och visas inte.  
Om procenttecken förekommer i texten behandlas de som en del av texten.  
Exempel: a^2+b^2=c^2%% Pythagoras 'sats  
Anvisningar för %PRODUCTNAME Math  
Mata in och redigera formler  
Mata in radbrytning  
Så här skriver du en formel på två rader i %PRODUCTNAME Math (med manuell radbrytning).  
En radbrytning uppnår man med kommandot "newline".  
Allt som står efter detta finns på en ny rad.  
Mata in parenteser  
Kan parenteser i %PRODUCTNAME Math även visas enskilt och i fritt definierbar storlek?  
Med "left" och "right "kan du visserligen sätta enskilda parenteser, men då har parenteserna ingen fast storlek eftersom de anpassar sig till argumentet.  
Men det finns en möjlighet att visa enskilda parenteser med fast storlek.  
Ett omvänt snedstreck "\" (backslash) sätts framför de normala parenteserna.  
De här parenteserna beter sig då som vilken annan symbol som helst och har inte längre den speciella funktionen för parenteser, d.v.s. de har inte en grupperande verkan och justeringen är som vid andra symboler, jfr. "left lbrace x right none" och "size *2 langle x rangle "och "size *2 \langle x \rangle".  
Om du vill pröva exemplen måste du mata in dem utan citationstecken.  
Välkommen till %PRODUCTNAME Math-hjälpen  
Hjälp till %PRODUCTNAME Math  
Referens  
Hjälp till hjälpen  
Menyer  
Menylisten innehåller alla kommandon som du behöver när du arbetar med %PRODUCTNAME Math.  
Via den når du en lista över tillgängliga operatorer och kommandon för redigering, visning, placering, formatering, utskrift etc. av formeldokument och objekt som de innehåller.  
De flesta menypunkterna är bara tillgängliga när du skapar eller redigerar en formel.  
Arkiv  
I den här menyn hittar du allmänna kommandon för hantering av formeldokument som t.ex. Öppna, Spara och Skriv ut.  
Öppna...  
AutoPilot  
I dessa dokument kan du sedan, om du vill, infoga sparade formler.  
Spara som...  
Versioner...  
Dokument som e-post...  
Egenskaper...  
Skriv ut...  
Skrivarinställning...  
Redigera  
Den innehåller dels allmänna kommandon, t.ex. för kopiering av innehåll, dels kommandon som är specifika för %PRODUCTNAME Math som t.ex. sökning efter platshållare eller stöd vid felsökning.  
Visa  
Här ställer du in visningsskalan och väljer vilka andra element som ska synas.  
De flesta kommandon som du kan ange i fönstret Kommandon kan du infoga genom att klicka med musen när du har öppnat urvalsfönstret med kommandot Visa - Urval.  
Skala  
Format  
Här hittar du kommandon som används till att formatera formler.  
Teckensnitt...  
Teckenstorlekar...  
Avstånd...  
Justering...  
Verktyg  
Här kan du öppna och redigera en symbolkatalog eller importera en extern formel som fil.  
Dessutom kan du ändra standardinställningarna för programmet här.  
Importera formel...  
Anpassa...  
Fönster  
Där finns även en lista över öppna dokument.  
Symbollister  
Här beskrivs symbollisterna som du kan använda när ett %PRODUCTNAME Math-dokument är öppet.  
Du kan anpassa alla lister efter dina behov, flytta eller radera ikoner eller infoga nya ikoner.  
Om du ändrar symbollisterna kommer naturligtvis konfigurationen att skilja sig mer eller mindre från den som beskrivs här.  
Statuslist  
På statuslisten visas information om det aktuella dokumentet.  
Du kan konfigurera den (under Verktyg - Anpassa...).  
Följande fält visas enligt standardinställningen:  
Verktygslist  
Verktygslisten innehåller viktiga funktioner som du ofta har användning av.  
Formelmarkör  
Funktioner i %PRODUCTNAME %PRODUCTVERSION Math  
Här får du en kort överblick över några viktiga funktioner i %PRODUCTNAME Math.  
De är överskådligt ordnade i ett urvalsfönster och du kan lätt infoga dem i ditt arbete genom att klicka på dem.  
Dessutom innehåller hjälpen en uttömmande referenslista och många användningsexempel.  
Skapa en formel  
Formler skapar du, precis som diagram och eventuellt även bilder, oftast inne i ett annat dokument.  
Om du fogar in en formel i ett annat dokument startas %PRODUCTNAME Math automatiskt.  
Du skapar, redigerar och formaterar formeln som du vill med hjälp av ett stort antal fördefinierade symboler och funktioner.  
Mata in en formel direkt  
Om du redan kan språket i %PRODUCTNAME Math, kan du även mata in en formel direkt.  
Markera sedan omskrivningen och välj motsvarande menypunkt. %PRODUCTNAME omvandlar då automatiskt den här texten till en formaterad formel.  
Det går inte att utvärdera eller beräkna formler här eftersom detta inte är ett kalkylprogram utan en formeleditor, d.v.s. en modul där du kan skriva och visa formler.  
Använd tabelldokument när du vill beräkna formler eller räknefunktionen i textdokument för lättare räkneuppgifter.  
Skapa en formel i kommandofönstret  
Du redigerar beskrivningen av formeln i kommandofönstret i %PRODUCTNAME Math.  
Formeln visas i textfönstret.  
Använd formelmarkören på verktygslisten för att inte tappa överblicken vid långa konstruktioner.  
I textfönstret visar den var du för tillfället befinner dig i kommandofönstret och omvänt.  
Om du klickar på ett ställe i något av fönstren markeras motsvarande plats i det andra fönstret.  
Individuella symboler  
Du kan skapa egna symboler och använda tecken från andra teckenuppsättningar.  
Till %PRODUCTNAME Maths baskatalog över tillgängliga tecken kan du lägga till ett valfritt antal nya och även sammanställa egna särskilda kataloger.  
Det finns många specialtecken (t.ex. halva klammerparenteser) som du kan använda.  
Använd snabbmenyerna  
Utnyttja möjligheterna som snabbmenyerna ger.  
Du öppnar dem med höger musknapp.  
Kommandofönstrets meny innehåller inte bara de kommandon som finns i urvalsfönstret utan även andra kommandon.  
Då slipper du att göra inmatningar i kommandofönstret via tangentbordet.  
Så hittar du den här funktionen...  
Textanpassning av  
Textanpassning på  
Textgenomflöde  
Hopp till föregående skript  
Hopp till nästa skript  
Menyn Arkiv  
Menyn Arkiv - Skicka - Disposition till presentation  
Menyn Arkiv - Skicka - Disposition till urklippet  
Menyn Arkiv - Skicka - Skapa AutoUtdrag  
Menyn Arkiv - Skicka - AutoUtdrag till presentation  
Menyn Arkiv - Skicka - Skapa HTML-dokument  
Menyn Arkiv - Skicka - Skapa HTML-dokument - Formatmall, menyn Arkiv - Skicka - Skapa samlingsdokument - Formatmall  
Menyn Arkiv - Kopplad utskrift..  
Ikon på databaslisten:  
Kopplad utskrift...  
Menyn Arkiv - Kopplad utskrift..., välj "E-post", klicka på... till höger om Bilagor.  
Menyn Redigera  
Menyn Redigera - AutoText...  
Kommando Ctrl +F3  
Ikon på verktygslisten:  
Redigera AutoText  
Menyn Redigera - Byt databas...  
Menyn Redigera - FÃ¤ltkommando...  
Menyn Redigera - Fotnot...  
Menyn Redigera - Förteckningspost...  
Snabbmenyn Förteckningspost...  
Menyn Format - OmrÃ¥den...  
Menyn Redigera - AutoText... - AutoText - Byt namn  
Menyn Redigera - LitteraturfÃ¶rteckningspost...  
Menyn Visa  
Menyn Visa - Linjal  
Menyn Visa - TextbegrÃ¤nsningar  
Menyn Visa - Markeringar  
Kommando Ctrl +F8  
Menyn Visa - Fältkommandon  
Tangentkombinationen Kommando Ctrl +F9  
Menyn Visa - Kontrolltecken  
Kommando Ctrl +F10  
Ikon på verktygslisten:  
Kontrolltecken på / av  
Menyn Visa - Onlinelayout  
Ikon på verktygslisten:  
Onlinelayout  
Menyn Visa - Utskriftslayout  
Ikon på verktygslisten / web:  
Utskriftslayout på / av  
Menyn Visa - Dolda stycken  
Menyn Infoga  
Menyn Infoga - Manuell brytning...  
Menyn Infoga - Fältkommando  
Snabbmenyn Fältkommando... (vid infogat fältkommando)  
Menyn Infoga - FÃ¤ltkommando - Datum  
Menyn Infoga - FÃ¤ltkommando - Klockslag  
Menyn Infoga - FÃ¤ltkommando - Sidnummer  
Menyn Infoga - FÃ¤ltkommando - Sidantal  
Menyn Infoga - FÃ¤ltkommando - Ã„mne  
Menyn Infoga - FÃ¤ltkommando - Titel  
Menyn Infoga - FÃ¤ltkommando - FÃ¶rfattare  
Menyn Infoga - Fältkommando - Andra...  
Dubbelklicka i det stora fältet till höger i statuslisten när inget är markerat  
Kommando Ctrl +F2  
Ikon på verktygslisten:  
Infoga fältkommandon  
Menyn Infoga - Fältkommando - Andra... - fliken Dokument  
Menyn Infoga - Fältkommando - Andra... - fliken Referenser  
Menyn Infoga - Korshänvisning  
Menyn Infoga - Fältkommando - Andra... - fliken Funktioner  
Menyn Infoga - Fältkommando - Andra... - fliken Dokumentinfo  
Menyn Infoga - Fältkommando - Andra... - fliken Variabler  
Menyn Infoga - Fältkommando - Andra... - fliken Databas  
Menyn Infoga - Område...  
Ikon på utrullningslisten Infoga på verktygslisten och på verktygslisten / web  
Infoga område  
Menyn Infoga - Område... - fliken Område och menyn Format - OmrÃ¥den...  
Fotnot: menyn Infoga - Fotnot...  
Snabbmenyn Fotnot... (vid infogad fot - / slutnot)  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga fotnot direkt  
Infoga slutnot direkt  
Menyn Infoga - Bildtext...  
Snabbmenyn Bildtext...  
Menyn Infoga - Bildtext... - Alternativ  
Snabbmenyn Bildtext... - Alternativ  
Menyn Infoga - Bokmärke...  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga bokmärke  
Menyn Infoga - Skript (bara vid HTML-dokument)  
Menyn Infoga - FÃ¶rteckningar  
Menyn Infoga - Förteckningar - Post...  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga indexmarkering  
Menyn Infoga - FÃ¶rteckningar - FÃ¶rteckningar...  
Menyn Infoga - FÃ¶rteckningar - LitteraturfÃ¶rteckningspost...  
Menyn Infoga - FÃ¶rteckningar - FÃ¶rteckningar...  
Menyn Infoga - Förteckningar - Förteckningar... - fliken FÃ¶rteckning  
Menyn Infoga - Förteckningar - Förteckningar... - fliken Förteckning (beroende på vald förteckningstyp)  
Menyn Infoga - Förteckningar - Förteckningar... - (fliken Förteckning när typen Innehållsförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... - (fliken Förteckning när typen Sakregister är vald)  
Menyn Infoga - Förteckningar - Förteckningar... - (fliken Förteckning när typen Illustrationsförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... - (fliken Förteckning när typen Tabellförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... - (fliken Förteckning när typen Användardefinierad är vald)  
Menyn Infoga - Förteckningar - Förteckningar... - (fliken Förteckning när typen Objektförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... - (fliken Förteckning när typen Litteraturförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... - markera fältet "Ytterligare mallar" och klicka sedan på...  
Menyn Infoga - Förteckningar - Förteckningar... fliken Poster (beroende på vald förteckningstyp)  
Menyn Infoga - Förteckningar - Förteckningar... (fliken Poster när typen Innehållsförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... (fliken Poster när typen Sakregister är vald)  
Menyn Infoga - Förteckningar - Förteckningar... (fliken Poster när typen Illustrationsförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... (fliken Poster när typen Tabellförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... (fliken Poster när typen Användardefinierad är vald)  
Menyn Infoga - Förteckningar - Förteckningar... (fliken Poster när typen Objektförteckning är vald)  
Menyn Infoga - Förteckningar - Förteckningar... (fliken Poster när typen Litteraturförteckning är vald)  
Menyn Infoga - Förteckningar - Litteraturförteckningspost... - kommandoknappen Redigera  
Menyn Infoga - Förteckningar - Förteckningar... - fliken Mallar  
Menyn Infoga - Kuvert...  
Menyn Infoga - Kuvert... - fliken Kuvert  
Menyn Infoga - Kuvert... - fliken Format  
Menyn Infoga - Kuvert... - fliken Skrivare  
Menyn Infoga - Ram...  
Menyn Format - Ram...  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga ram manuellt  
Menyn Infoga - Tabell...  
Kommando Ctrl +F12  
Ikon på utrullningslisten Infoga på verktygslisten:  
Infoga tabell  
Menyn Infoga - Horisontell linje...  
Menyn Infoga - Fil...  
Ikon på utrullningslisten Infoga på verktygslisten:  
Dokument  
Menyn Infoga - Sidhuvud  
Menyn Infoga - Sidfot  
Menyn Format  
Menyn Format - Stycke... - fliken AnfangsbokstÃ¤ver  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken AnfangsbokstÃ¤ver  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken AnfangsbokstÃ¤ver  
Menyn Format - Stycke... - fliken TextflÃ¶de  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken TextflÃ¶de  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken TextflÃ¶de  
Menyn Redigera - Sök och ersätt... - Format... - fliken TextflÃ¶de  
Menyn Format - Sida...  
Menyn Format - Mallar - Katalog... - Nytt... / Ändra... (vid sidformatmallar)  
Menyn Format - Stylist - snabbmenyn Nytt... / Ändra... (vid sidformatmallar)  
Menyn Format - Stycke... - fliken Numrering  
Menyn Format - Mallar - Katalog... - Nytt... / Ändra... (vid styckeformatmallar) - fliken Numrering  
Menyn Format - Stylist - snabbmenyn Nytt... / Ändra... (vid styckeformatmallar) - fliken Numrering  
Menyn Format - Områden... - kommandoknappen Alternativ  
Menyn Format - Sida... - fliken Kolumner  
Menyn Format - Ram... - fliken Kolumner  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Kolumner  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Kolumner  
Menyn Infoga - Ram... - fliken Kolumner  
Menyn Infoga eller Format - Områden... - fliken Kolumner  
Menyn Format - Sida... - fliken Fotnot  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Fotnot  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Fotnot  
Menyn Infoga - Område... - fliken Fot - / slutnoter  
Menyn Format - Områden... - kommandoknappen Alternativ - fliken Fot - / slutnoter  
Menyn Format - Mallar - Ladda...  
Menyn Format - Mallar - Katalog... - Nytt... / Ändra... (vid styckeformatmallar)  
Menyn Format - Stylist - snabbmenyn Nytt... / Ändra... (vid styckeformatmallar)  
Menyn Format - Mallar - Katalog... - Nytt... / Ändra... (vid teckenformatmallar)  
Menyn Format - Stylist - snabbmenyn Nytt... / Ändra... (vid teckenformatmallar)  
Menyn Format - Mallar - Katalog... - Nytt... / Ändra... (vid ramformatmallar)  
Menyn Format - Stylist - snabbmenyn Nytt... / Ändra... (vid ramformatmallar)  
Menyn Format - Mallar - Katalog... - Nytt... / Ändra... (vid numreringsformatmallar)  
Menyn Format - Stylist - snabbmenyn Nytt... / Ändra... (vid numreringsformatmallar)  
Menyn Format - Mallar - Katalog... - Nytt... (vid styckeformatmallar) - fliken Villkor  
Menyn Format - AutoFormat - Under inmatningen  
Menyn Format - AutoFormat  
Menyn Format - AutoFormat - AnvÃ¤nd  
Menyn Format - AutoFormat - AnvÃ¤nd och redigera Ã¤ndringar  
Meny Format - AutoFormat... (med markören i en tabell)  
Menyn Format - Grafik...  
Menyn Infoga - Grafik - Från fil... - Egenskaper  
Menyn Infoga - Grafik - Från fil... (när en grafik är markerad)  
Ikon på objektlisten (vid markerad grafik):  
Grafikegenskaper  
Menyn Format - Grafik... - fliken Typ  
Menyn Format - Objekt... - fliken Typ  
Menyn Format - Ram - fliken Typ  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Typ  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Typ  
Menyn Infoga - Ram... - fliken Typ  
Menyn Format - Grafik... - fliken Textanpassning  
Menyn Format - Objekt... - fliken Textanpassning  
Menyn Format - Ram... - fliken Textanpassning  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken Textanpassning  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken Textanpassning  
Menyn Infoga - Ram... - fliken Textanpassning  
Menyn Format - Textanpassning  
Menyn Format - Textanpassning - Redigera kontur...  
Menyn Format - Grafik... - fliken HyperlÃ¤nk  
Menyn Format - Ram... - fliken HyperlÃ¤nk  
Menyn Format - Objekt... - fliken HyperlÃ¤nk  
Menyn Infoga - Ram... - fliken HyperlÃ¤nk  
Menyn Format - Grafik... - fliken TillÃ¤gg  
Menyn Format - Objekt... - fliken TillÃ¤gg  
Menyn Format - Ram... - fliken TillÃ¤gg  
Menyn Format - Mallar - Katalog... - Ändra / Nytt... - fliken TillÃ¤gg  
Menyn Format - Stylist - snabbmenyn Ändra / Nytt... - fliken TillÃ¤gg  
Menyn Infoga - Ram... - fliken TillÃ¤gg  
Menyn Format - Grafik... - fliken Grafik  
Menyn Infoga / Format - Grafik... - fliken Makro  
Menyn Infoga / Format - Ram... - fliken Makro  
Menyn Format - Objekt... - fliken Makro  
Menyn Redigera - AutoText... - AutoText - Makro...  
Menyn Redigera - Image map - snabbmenyn - Makro...  
Menyn Infoga - Hyperlänk - kommandoknappen Händelser...  
Menyn Format - Tecken... - fliken Hyperlänk - Händelser...  
Menyn Format - Tabell...  
Menyn Format - Dela tabell...  
Menyn Format - Förbind tabeller  
Menyn Format - Tabell... - fliken Tabell  
Menyn Format - Tabell... - fliken Kolumner  
Menyn Format - Tabell... - fliken Textflöde  
Menyn Format - Cell  
Menyn Format - Cell - Förbinda  
Ikon på objektlisten:  
Förbind celler  
Menyn Format - Cell - Dela...  
Ikon på objektlisten:  
Dela cell  
Menyn Format - Cell - Skydda  
Menyn Format - Cell - Upphäv skydd  
Snabbmenyn i Navigator för tabeller  
Menyn Format - Cell - Överst  
Menyn Format - Cell - Mitten  
Menyn Format - Cell - Underst  
Menyn Format - Rad  
Menyn Format - Rad - Höjd...  
Menyn Format - Rad - Optimal höjd  
Ikon på utrullningslisten Optimera på objektlisten:  
Optimal radhöjd  
Menyn Format - Rad - Fördela jämnt  
Ikon på utrullningslisten Optimera på objektlisten:  
Fördela raderna jämnt  
Menyn Format - Rad - Välj ut  
Menyn Format - Rad - Radera  
Ikon på objektlisten:  
Radera rad  
Menyn Format - Kolumn  
Menyn Format - Kolumn - Bredd...  
Menyn Format - Kolumn - Optimal bredd  
Ikon på utrullningslisten Optimera på objektlisten:  
Dubbelklicka på den högra kolumnavgränsaren i kolumnhuvudena  
Optimal kolumnbredd  
Menyn Format - Kolumn - Fördela jämnt  
Ikon på utrullningslisten Optimera på objektlisten:  
Fördela kolumnerna jämnt  
Menyn Format - Kolumn - Välj ut  
Menyn Format - Kolumn - Infoga...  
Menyn Format - Rad - Infoga...  
Ikon på objektlisten:  
Infoga kolumn  
Infoga rad  
Menyn Format - Kolumn - Radera  
Ikon på objektlisten:  
Radera kolumn  
Menyn Format - Objekt...  
Ikon på objektlisten (när ett objekt är markerat):  
Objektegenskaper  
Ramegenskaper  
Menyn Verktyg  
Menyn Verktyg - Avstavning...  
Menyn Verktyg - Kapitelnumrering...  
Menyn Verktyg - Kapitelnumrering... fliken Numrering  
Menyn Verktyg - Radnumrering...  
Menyn Verktyg - Fotnoter...  
Menyn Verktyg - Fotnoter... fliken Fotnoter  
Menyn Verktyg - Fotnoter... fliken Slutnoter  
Menyn Verktyg - Text <-> Tabell...  
Menyn Verktyg - Sortera...  
Menyn Verktyg - Beräkna  
Tangentkombinationen Kommando Ctrl +plustecken  
Menyn Verktyg - Uppdatera  
Menyn Verktyg - Uppdatera - Sidformatering  
Menyn Verktyg - Uppdatera - Aktuell fÃ¶rteckning  
Menyn Verktyg - Uppdatera - Alla fÃ¶rteckningar  
Menyn Verktyg - Uppdatera - Uppdatera allt  
Menyn Verktyg - Uppdatera - Fält  
Tangenten F9  
Menyn Verktyg - Uppdatera - LÃ¤nkar  
Menyn Verktyg - Uppdatera - Alla diagram  
Kopplad utskrift  
Här hittar du alla funktioner för att skriva ut och spara standardbrev.  
Innan du använder det här kommandot väljer du den länkade datakällan varifrån t.ex. adresser ska hämtas och infogas i motsvarande fält i dokumentet.  
Själva utskriften startar du i dialogrutan Kopplad utskrift.  
Databasinformationen infogas först vid utskriften vid databasfältkommandonas (platshållarnas) positioner.  
Information om att infoga databasfältkommandon finns under Infoga - Fältkommando - Andra under fliken Databas.  
Dataposter  
Här anger du antalet dataposter för den kopplade utskriften.  
Ett brev skrivs ut för varje datapost.  
Alla  
Alla dataposter i databasen (databasfrågan) behandlas.  
Markerade dataposter  
Det här alternativfältet kan du bara välja om du tidigare har markerat motsvarande dataposter i databasen.  
Från:  
Här väljer du vilka dataposter som ska tas med i den kopplade utskriften.  
Från:  
Här anger du numret på den första dataposten som ska användas vid utskriften.  
Till:  
Här anger du numret på den sista dataposten som ska användas vid utskriften.  
Utdata  
Här väljer du om den kopplade utskriften ska göras direkt, om du ska skicka den elektroniskt via e-post till mottagarnas adresser i adressboken eller om du först vill skapa en fil av den.  
Skrivare  
Välj det här alternativet om standardbreven ska skrivas ut.  
E-post  
Välj det här alternativet om standardbreven ska skickas med e-post.  
Du kan då välja uppgifter i Adressfält et och i textfältet Angående samt ange e-postformatet under E-postformat.  
Fil  
Markera det här alternativet om du vill göra en fil av den kopplade utskriften.  
Skapa enstaka utskriftsjobb  
I annat fall skickas standardbreven som ett enda utskriftsjobb.  
Adressfält  
Här väljer du det datafält i databasen där e-postadressen finns.  
Angående  
Här anger du ärenderubriken.  
Bilagor  
Filnamnen är åtskiljda av semikolon.  
Med kommandoknappen... kan du öppna dialogrutan Välj ut filer där du kan välja filerna som ska bifogas.  
E-postformat  
Här anger du med vilket e-postformat den kopplade utskriften ska skapas.  
%PRODUCTNAME Writer  
Om du markerar den här kryssrutan, skapas den kopplade utskriften förutom i ASCII-format även i %PRODUCTNAME Writer-format.  
HTML  
Om du klickar i den här kryssrutan, ger du dessutom den kopplade utskriften HTML -format.  
RTF  
Klicka här om du vill att även RTF -format ska användas.  
Sökväg  
Här anger du den katalog där filen med den kopplade utskriften ska skapas.  
...  
Med den här kommandoknappen öppnar du en dialogruta där du kan välja mapp.  
Generera filnamn från - Databasfält  
Markera det här alternativet om innehållet i de markerade datafälten ska användas som filnamn.  
Generera filnamn från - Anpassa  
Markera det här alternativet om filnamnen ska skapas på basis av den text som du skriver i textfältet samt löpnummer.  
Välj ut filer  
Här markerar du de filer du vill bifoga.  
Filer  
Här visas de filer som lagts till i den här dialogrutan.  
Lägg till...  
Om du klickar på Lägg till, kan du i dialogrutan Öppna markera en fil som läggs till i fillistan.  
Radera  
Klicka på Radera, om du vill ta bort den markerade filen från listan.  
Disposition till presentation  
Med det här kommandot överför du det aktuella dokumentets disposition till ett nytt presentationsdokument.  
Disposition till urklipp  
Med det här kommandot kopierar du dispositionen för det aktuella dokumentet till urklippet i Rich Text Format (RTF).  
Skapa AutoUtdrag  
Här kopierar du överskrifterna och ett antal följande stycken i det aktuella dokumentet till ett nytt AutoUtdrag-textdokument.  
AutoUtdrag ger bättre överblick över långa dokument.  
Du kan ställa in antalet kapitelnivåer och antalet stycken som ska visas per kapitelnivå.  
Alla nivåer och stycken som ligger under respektive inställning döljs.  
Inkluderade kapitelnivåer  
Här anger du antalet steg för nivåerna som ska kopieras till det nya dokumentet.  
Om du t.ex. väljer 4 nivåer, så övertas de stycken som är formaterade med överskrift 1 till överskrift 4, och efter varje stycke övertas det antal följande stycken som du har angett i fältet Stycken per kapitel.  
Stycken per kapitel  
Med de här rotationsknapparna definierar du det maximala antalet på varandra följande stycken som ska övertas till AutoUtdrag-textdokumentet efter varje inkluderad överskrift.  
Av det angivna antalet övertas högst så många stycken som krävs för att nå nästa stycke med formateringen "Överskrift".  
AutoUtdrag till presentation  
Med det här kommandot överför du ett AutoUtdrag som disposition till ett nytt presentationsdokument.  
AutoUtdrag hjälper dig att ge långa dokument en överskådlig utformning.  
Inkluderade kapitelnivåer  
Här anger du antalet steg för de nivåer som ska kopieras till det nya dokumentet.  
Efter varje stycke överförs det antal efterföljande stycken som du har angett i fältet Stycken per kapitel.  
Stycken per kapitel  
Med de här rotationsknapparna definierar du det maximala antalet på varandra följande stycken som ska överföras till AutoUtdrag-textdokumentet efter varje inkluderad överskrift.  
Av det angivna antalet överförs högst så många stycken som krävs för att nå nästa stycke med formateringen "Överskrift".  
HTML-dokumentets namn och sökväg  
Om du väljer Arkiv - Skicka - Skapa HTML-dokument delas det aktuella dokumentet upp i en rad HTML-dokument som är ihopkopplade med hyperlänkar.  
Dokumenten delas vid de stycken som är formaterade med en viss formatmall.  
En fildialogruta visas, där du anger katalog och namn för huvuddokumentet som ska skapas.  
Deldokumenten får automatiskt namn, som består av huvuddokumentets namn och ett löpnummer.  
Titeln på en nyskapad fil tas automatiskt upp i dokumentinformationen.  
Den hämtas från eventuellt befintlig titel och från kapitelöverskriften.  
Visningsområde  
Filnamn  
Aktuell formatmall  
Välj styckeformatet som ska fungera som avgränsning.  
I normala fall delar du utgångsdokumentet vid de stycken som har formaterats med formatet "Överskrift 1".  
På så vis blir varje kapitel till ett eget deldokument.  
Här kan du också välja en annan mall bland styckeformatmallarna som används i dokumentet.  
Filtyp  
Spara  
Automatiskt filnamnstillägg  
Navigator  
Med den här funktionen sätter du på och stänger av Navigator.  
Med den tar du dig snabbt till särskilda kapitel och objekt, och du kan bl.a. ordna kapitel och infoga objekt från andra öppna dokument.  
På snabbmenyn till posterna i Navigator visas särskilda kommandon, t.ex. för att redigera, byta namn, upphäva tabellskydd, omvandla en innehållsförteckning till normal text och mycket annat.  
Navigator är ett förankringsbart fönster.  
När Du vill att Navigator ska visas på bildskärmen och Du har ett dokument öppet väljer Du Redigera - Navigator, klickar på ikonen på funktionslisten eller trycker på F5.  
Om Navigator täcker viktiga textpartier, kan Du flytta fönstret genom att peka på rubrikraden, trycka ned vänster musknapp och dra.  
Om Du vill förankra Navigator mot fönsterkanten, håller Du Kommando Ctrl -tangenten nedtryckt när Du flyttar.  
Du kan förankra och frigöra Navigator direkt genom att trycka på Kommando Ctrl-tangenten och dubbelklicka i ett fritt område i Navigator-fönstret.  
I Navigator förtecknas olika element som kan finnas i dokumenten.  
Om det aktuella dokumentet innehåller element av en viss typ, visas detta i Navigator med ett litet plustecken framför motsvarande post.  
Om Du låter muspekaren stanna ett ögonblick på en sådan post, visar tipshjälpen - (menykommando Hjälp - Tips) hur många element av den här typen i som finns dokumentet.  
Om Du klickar på plustecknet framför en post, visas en lista över vilka element som finns i dokumentet.  
Om Du dubbelklickar på ett sådant element flyttas markören till motsvarande plats i dokumentet.  
Om ett dokumentinnehåll finns i dolda områden, visas bara det här innehållet i grått i Navigator.  
Tipshjälpen visar den dolda texten.  
Samma sak gäller för innehåll som finns i sidhuvuden eller sidfötter i sidformatmallar som inte används.  
Du kan hitta dolt innehåll, om det finns något, under tabeller, textramar, grafik, OLE-objekt, områden och förteckningar i Navigator.  
Om Du vill ändra ett visst element i dokumentet, öppnar Du bara snabbmenyn till motsvarande element i Navigator och väljer kommandot Redigera....  
Kommandot öppnar dialogrutan för respektive element, så att Du kan redigera det.  
För tabeller kan du dessutom upphäva ett aktiverat cellskydd.  
Om du har skyddat en eller flera celler med kommandot Format - Cell - Skydda så att de inte kan redigeras, kan du ta bort detta skydd via tabellpostens snabbmeny, där Du väljer Tabell - Upphäv skydd.  
Med kommandot Upphäv förteckning på en förtecknings snabbmeny gör du t.ex. om en innehållsförteckning till normal text.  
Med kommandot Skrivskyddad, som kan vara bockmarkerat, aktiverar och inaktiverar Du skrivskyddet för t ex en förteckning.  
Med kommandot Radera på ett markerat objekts snabbmeny raderar Du objektet från dokumentet.  
Du kan även använda tangenten Delete.  
Med kommandot Byt namn på ett markerat objekts snabbmeny i Navigator öppnar Du en dialogruta där Du kan ge objektet ett nytt namn.  
Om Du snabbt vill komma till en viss innehållstyp i dokumentet kan Du även använda utrullningslisten Navigation, som Du öppnar genom att klicka på ikonen Navigation.  
Denna ikon finns både i Navigator och nedtill på höger bildrullningslist i ett öppet textdokument.  
Växla  
Med den här ikonen växlar du mellan samlingsläge och normalläge.  
Den är bara aktiv om du har öppnat ett samlingsdokument (t.ex. med menykommandot Arkiv - Nytt - Samlingsdokument).  
Växla  
Navigation  
Genom att klicka på "Föregående objekt" och "Nästa objekt "kan Du bläddra mellan dem.  
Med utrullningslisten Navigation kan Du, förutom att välja objekttyp, också aktivera funktionen Fortsätta en sökning.  
Navigation  
Föregående objekt  
Med den här symbolen flyttar Du markören till nästa objekt i riktning mot dokumentets början.  
Det objekt dit Du vill komma kan Du ange på utrullningslisten Navigation.  
Namnet på ikonen beror av det valda objektets typ.  
Om Du med navigationssymbolen t ex väljer textramar, heter ikonen "Föregående textram".  
Föregående objekt  
Nästa objekt  
Med den här symbolen flyttar Du markören till nästa objekt i riktning mot dokumentets slut.  
Det objekt dit Du vill komma kan Du ange på utrullningslisten Navigation.  
Namnet på ikonen beror av det valda objektets typ.  
Om Du med navigationssymbolen t ex väljer textramar, heter ikonen "Nästa textram".  
Nästa objekt  
Sidnummer  
I det här rotationsfältet kan Du ange ett sidnummer och bekräfta det med returtangenten.  
Markören flyttas till början av den valda sidan.  
Med tangenterna PageUp (PgUp) och PageDown (PgDn) anger Du i rotationsfältet numret på den sista och den första sidan.  
Sidnumret är markerat, så att du direkt kan skriva det nya sidnumret och bekräfta det med returtangenten.  
Om Du ändrar numret i inmatningsfältet, flyttas markören i texten efter en liten fördröjning till den nya sidan.  
Sida  
Urvalsbox  
Med den här ikonen växlar Du mellan att visa och dölja det nedre Navigatorområdet, såvida Navigatorfönstret inte är förankrat.  
Urvalsbox på / av  
Växla innehållsvisning  
Med den här ikonen växlar Du i Navigator mellan att visa alla element eller bara de element som är markerade i Navigator med den aktuella markören.  
Växla innehållsvisning  
Det är bara om den här ikonen är intryckt som du kan flytta överskrifterna genom att dra och släppa dem i Navigator.  
På så vis flyttar du samtidigt motsvarande kapitel i dokumentet.  
Sätt temporärt bokmärke  
Med det här alternativet infogar Du ett temporärt bokmärke utan namn där markören står.  
Välj posten Temporärt bokmärke på utrullningslisten Navigation och gå sedan till bokmärkena med kommandoknapparna Nästa temporära bokmärke och Föregående temporära bokmärke.  
Sätt temporärt bokmärke  
Du kan infoga upp till fem temporära bokmärken samtidigt.  
Om Du infogar fler raderas det äldsta.  
Sidhuvud  
Med den här symbolen flyttar Du markören till sidhuvudet eller från sidhuvudet till dokumentets textområde.  
Sidhuvud  
Sidfot  
Med den här symbolen flyttar Du markören fram och tillbaka mellan sidfoten och dokumentets textområde.  
Sidfot  
Ankare <-> Text  
Med den här symbolen flyttar Du markören fram och tillbaka mellan fotnotsområdet och fotnotsmärket.  
Ankare <-> Text  
Draläge  
Om du klickar på den här ikonen visas en undermeny där du kan välja draläge.  
Du kan även öppna undermenyn via snabbmenyn på Navigators visningsområde.  
Här bestämmer du vilken åtgärd som ska utföras när du drar och släpper ett element från Navigator till ett dokument.  
Ikonen byter utseende alltefter draläget och visar på det viset direkt om en hyperlänk, en länk eller en kopia kommer att skapas.  
Draläge  
Infoga som hyperlänk  
Om Du har markerat den här posten, skapas en hyperlänk när Du drar ett objekt till ett %PRODUCTNAME -dokument.  
Du kan klicka på den här hyperlänken om Du vill hoppa till det element vars symbol Du just har skapat med dra-och-släpp.  
Infoga som länk  
Om Du har markerat den här posten, skapas en länk när Du drar ett objekt till ett %PRODUCTNAME -dokument.  
I ett %PRODUCTNAME -textdokument skapas elementet som skyddat område.  
Om elementet i källdokumentet ändras, ändras också innehållet i det länkade området nästa gång Du öppnar måldokumentet eller när Du uppdaterar innehållet i det länkade området i dialogrutan Redigera - Länkar...  
Det går inte att länka grafikobjekt, OLE-objekt, referenser eller förteckningar.  
Infoga som kopia  
Om Du har markerat den här posten, innebär det att om Du drar och släpper ett element till ett %PRODUCTNAME -dokument, skapas en kopia av elementet.  
Det blir då ett icke skyddat område.  
Det går inte att kopiera grafikobjekt, OLE-objekt, referenser eller förteckningar.  
Visade överskriftsnivåer  
Om Du klickar på den här ikonen öppnas en undermeny, där Du kan välja vilka överskriftsnivåer som ska visas.  
Den här undermenyn kan Du också öppna via snabbmenyn i Navigators visningsområde under Dispositionsnivåer.  
1-10  
Om Du väljer 10, visas alla tio nivåerna.  
Visade överskriftsnivåer  
Kapitel uppåt  
Det kapitel som är markerat i Navigator-fönstret förflyttas - tillsammans med tillhörande underkapitel - ett steg i riktning mot dokumentets början.  
Om Du vill flytta enbart det markerade kapitlet, håller Du Kommando Ctrl -tangenten nedtryckt samtidigt som Du klickar på ikonen.  
Kapitel uppåt  
Kapitel nedåt  
Det kapitel som är markerat i Navigator-fönstret förflyttas - tillsammans med tillhörande underkapitel - ett steg i riktning mot dokumentets slut.  
Om Du vill flytta enbart det markerade kapitlet, håller Du Kommando Ctrl -tangenten nedtryckt samtidigt som Du klickar på ikonen.  
Kapitel nedåt  
När Du vidtar den här åtgärden flyttas även texten mellan kapitelrubrikerna.  
Höj nivån  
Den kapitelrubrik som är markerad i Navigator-fönstret flyttas - tillsammans med tillhörande undernivåer - en nivå uppåt.  
Om Du vill flytta enbart det markerade kapitlet, håller Du Kommando Ctrl -tangenten nedtryckt samtidigt som Du klickar på ikonen.  
Höj nivån  
Sänk nivån  
Den kapitelrubrik som är markerad i Navigator-fönstret flyttas - tillsammans med tillhörande undernivåer - en nivå nedåt.  
Om Du vill flytta enbart det markerade kapitlet, håller Du Kommando Ctrl -tangenten nedtryckt samtidigt som Du klickar på ikonen.  
Sänk nivån  
Laddade dokument  
I den här listrutan nedtill i Navigator visas namnen på de laddade dokumenten.  
Om Du vill byta till visning av uppgifter i ett annat laddat dokument, klickar Du på dokumentnamnet.  
Efter varje dokumentnamn visas inom parentes om det är aktivt eller inaktivt.  
Det aktiva dokumentet väljer Du på menyn Fönster.  
På Navigatorfönstrets snabbmeny finns kommandot Visa, med vilket du öppnar en undermeny som innehåller samma alternativ som listrutan Laddade dokument.  
Här väljer du vilket dokument som Navigator ska visa information om.  
Om du väljer posten Aktivt fönster, ändras visningen i Navigator automatiskt om du byter aktuellt dokument.  
Navigation  
Om du klickar på den här ikonen i Navigator eller nere till höger vid dokumentfönstrets kant, öppnas en utrullningslist där du kan välja bland målen som finns i dokumentet.  
Sedan kan du flytta textmarkören till föregående eller nästa mål i dokumentet genom att trycka på pilknapparna som finns direkt ovanför och nedanför ikonen.  
Så länge Du inte har valt någon annan post, hoppar Du, enligt standardinställningen, med pilknapparna till föregående eller nästa sida i dokumentet.  
De båda dubbelpil-symbolerna är svarta om Du bläddrar igenom sidor, och blå om Du hoppar till andra objekt.  
Posterna överensstämmer i stor utsträckning med dem i Navigator -rutan.  
Dessutom kan Du även välja andra hoppadresser, t ex temporära bokmärken som Du kan sätta med ikonen Sätt temporärt bokmärke i Navigator.  
I utrullningslisten Navigation kan Du välja något av följande alternativ som objekt: tabell, textramar, grafik, OLE-objekt, sida, överskrift, temporärt bokmärke, ritobjekt, kontrollfält, område, bokmärke, markering, fotnot, anteckning, förteckningspost eller (felaktig) tabellformel.  
När det gäller tabellformler kan Du antingen hoppa till alla tabellformler som finns i dokumentet eller bara till de felaktiga.  
Formler med följdfel (alltså sådana som refererar till felaktiga formler) ignoreras.  
Så här arbetar Du med utrullningslisten Navigation  
Öppna utrullningslisten Navigation genom att klicka på ikonen längst ned på bildrullningslisten.  
Om Du behöver använda utrullningslisten ofta, och om det finns gott om plats på bildskärmen, kan Du flytta den från dess vanliga plats genom att dra den och placera den någon annanstans på skärmen.  
Klicka på ikonen för den typ av objekt som Du vill bläddra igenom.  
Pilknapparnas namn ändras beroende på vilken typ av objekt som Du har valt.  
Textmarkören flyttas då till det valda objektet.  
Välj menykommandot Verktyg - Anpassa.  
På de olika flikarna för anpassning av menyer, tangentbordskommandon och symbollister hittar Du olika funktioner för navigation inom dokumentet under kategorin "Navigera".  
Med funktionerna "Till nästa / föregående indexmarkering" kan Du t ex hoppa till förteckningsmarkeringarna i dokumentet.  
Upprepa sökning  
Med ikonen Upprepa sökning på utrullningslisten Navigation kan Du fortsätta en sökning som Du har startat via dialogrutan Sök och ersätt.  
Aktivera den fortsatta sökningen genom att klicka på ikonen.  
De blå pilknapparna på den vertikala bildrullningslisten får nu funktionerna Sök vidare framåt och Sök vidare bakåt.  
Om Du klickar på någon av pilknapparna, fortsätter sökningen efter det begrepp som Du har angett i dialogrutan Sök och ersätt.  
Observera att den här funktionen endast är tillgänglig om Du redan har genomfört en sökning.  
AutoText  
Med AutoText är det lätt att administrera textblock som innehåller texter som man ofta behöver, även med formatering, grafik, ramar och så vidare.  
Sedan kan du infoga textblock i ett dokument genom att ange deras tilldelade förkortning och trycka på funktionstangenten F3.  
Du kommer snabbt åt AutoTexter genom att klicka på ikonen Redigera AutoText på verktygslisten och hålla musknappen nedtryckt.  
Här visas AutoTexternas förkortningar och namn.  
AutoText  
Här visas de områden som Du har tillgång till samt namnen på de enskilda textblocken med tillhörande förkortningar.  
Tipshjälpen visar den fullständiga sökvägen och namnet för AutoText-områdena.  
Visa resten av namnet som tips vid inmatningen  
Om den här rutan är markerad, visas en tipshjälp när du matar in en ny text om de första tre tecken överensstämmer med namnet på ett AutoText-block.  
I tipshjälpen visas namnet på AutoText-blocket.  
Om du nu trycker på Retur, ersätts de inskrivna tecknen av motsvarande AutoText.  
När det gäller exemplet med blindtexten räcker det alltså att skriva Bli.  
I tipshjälpen visas då Blindtext, och när du trycker på Retur infogas blindtexten.  
Om det finns flera poster vars namn börjar med samma bokstäver, kan Du få fram även dem i tipshjälpen med kortkommandot Kommando Ctrl +tabbtangenten.  
Du bläddrar bakåt till redan visade poster med kortkommandot Kommando Ctrl +Skift+tabbtangenten.  
Namn  
Här visas en förteckning över alla namn på de textblock som är tillgängliga i detta område.  
Välj det namn Du vill ha.  
Förkortning  
I det här fältet visas bokstavskombinationen för det aktuella textblocket.  
Listruta  
Du får en bättre överblick om Du ordnar in varje textblock i ett område.  
I listrutan nedanför inmatningsfältet väljer Du önskat område.  
Fälten visas enligt samma mönster som i Explorer.  
Om Du klickar på symbolen visas allt innehåll, dvs alla tillhörande textblock.  
Om Du väljer ett av dem, visas det i inmatningsfältet.  
Genom att klicka på kommandoknappen Infoga eller dubbelklicka på en post för Du in det valda textblocket i dokumentet.  
Med musen kan Du enkelt dra och släppa textblock mellan områden.  
Infoga  
Om Du klickar på den här kommandoknappen, infogas det markerade textblocket i dokumentet där markören står.  
Du kan även infoga ett textblock utan att öppna menyn.  
Då skriver Du bara förkortningen och trycker på F3.  
När Du infogar oformaterade textblock övertas den styckeformatering som gäller för det stycke som Du infogar blocket i.  
AutoText  
Med det menykommando som visas när Du klickar på den här kommandoknappen kan Du utföra alla administrativa uppgifter.  
Nytt  
Den text som är markerad i dokumentet sparas i den aktuella textblocksfilen under den beteckning som är införd i fältet Namn.  
Det kommandot går bara att använda om Du har ändrat det som står under Namn och angett ett nytt namn.  
Ny (bara text)  
Den markerade texten infogas i AutoTexten på samma sätt som med Nytt.  
Eventuella formateringar, grafiska objekt, tabeller osv inkluderas inte.  
Kopiera  
Funktionen är särskilt intressant när det gäller längre textblock.  
Ersätt  
Innehållet i det textblock som är markerat under Namn ersätts med den text som är markerad i dokumentet.  
Byt namn  
Välj det här menykommandot om Du vill ändra den aktuella beteckningen på textblocket och / eller bokstavskombinationen i förkortningen.  
Det nya namnet anger Du i dialogrutan Byt namn på textblock.  
Redigera  
Innehållet i det textblock som är markerat under Namn visas i arbetsområdet och kan redigeras där.  
När Du har redigerat textblocket väljer Du Arkiv - Spara textblock och därefter Arkiv - Stäng.  
Makro...  
Med det här menykommandot öppnar Du dialogrutan Tilldela makro, där Du kan tilldela det aktuella textelementet körningen av ett makro.  
De makron som är kopplade till några av de AutoTexter som medföljer programmet kan Du använda för Dina egna AutoTexter.  
I de AutoTexter, som Du har sparat med alternativet "Enbart text", kan Du t ex infoga textsträngar som <field:company> eller <placeholder :"Text" :"Hjälptext ">.  
Makrona byter ut teckensträngarna mot motsvarande fältkommandon.  
Importera  
Då öppnas en dialogruta där du kan välja ett MS Word 97 / 2000-dokument eller en mall.  
Alla textblock som eventuellt finns i dem importeras som %PRODUCTNAME Writer AutoText-block.  
Områden...  
Om du vill få en bättre överblick kan du tilldela varje textblock ett område.  
Med den här kommandoknappen öppnar du dialogrutan Redigera områden.  
Redigera områden  
Här skapar du ett nytt område för textblock, döper om ett befintligt område eller raderar det.  
Område  
Ange här ett namn på ett nytt område eller ett område som ska ändras.  
Förutom alla bokstäver i alfabetet kan Du använda alla andra tecken som kan tas emot av filsystemet, vilket kan innebära att skillnad görs mellan versaler och gemener.  
I visningsfönstret visas det befintliga namnet.  
Genom att klicka på kommandoknappen Nytt skapar Du ett nytt område, och genom att klicka på kommandoknappen Byt namn kan Du ändra på namnet på ett befintligt område.  
Sökväg  
I det här fältet visas den aktuella sökvägen där AutoText-blocken är sparade.  
Välj här sökvägen där du vill spara din AutoText.  
Nytt  
När Du har skrivit ett nytt namn, kan Du använda den här kommandoknappen.  
Klicka på Nytt om Du vill införa det nya AutoText-området under det nya namnet.  
Byt namn  
Om Du skriver ett namn i inmatningsfältet Område får Du förutom kommandoknappen Nytt också tillgång till funktionen Byt namn.  
Klicka på den när ändringen ska införas.  
Tänk också på att stänga dialogrutan Redigera områden med knappen OK, så att alla redigeringar sparas.  
Urvalslista  
I fönstret visas de redan definierade områdena med tillhörande sökväg.  
När Du har infogat eller ändrat ett område visas även resultatet av de åtgärderna här.  
Detsamma gäller för radering av ett område.  
Sökväg...  
Med den här kommandoknappen öppnar Du dialogrutan Välj sökvägar.  
Om du vill använda fler sökvägar än standardsökvägen till AutoText, måste du lägga till dem under Sökväg... i dialogrutan AutoText eller under posten AutoText under Verktyg - Alternativ - %PRODUCTNAME - Sökvägar.  
Spara länkar relativt  
Du kan spara de länkar som finns i textblocket absolut (med angivande av lagringsenhet) eller relativt (dvs utgående från den mapp som innehåller AutoText-komponenterna).  
Att spara relativt kan vara praktiskt, t ex om Du sparar AutoTexter som är gemensamma för alla medarbetare på en nätverksserver, vilken kan mappas under olika enhetsbokstäver.  
I filsystemet  
Markera den här kryssrutan om Du vill att länkar till filer på Din egen dator ska anges med relativa adresser.  
På Internet  
Markera den här kryssrutan, om Du vill att länkar till filer på Internet (hyperlänkar) ska anges med relativa adresser.  
Visa förhandsvisning  
Med den här kryssrutan aktiverar och inaktiverar Du förhandsvisningen.  
Förhandsvisning  
I den här rutan visas en förhandsvisning av den valda AutoTexten.  
Byt namn på textblock  
Med den här dialogrutan kan Du byta namn på ett textblock som Du tidigare har markerat i dialogrutan AutoText.  
Namn  
I det här textfältet står namnet på det textblock som Du vill ändra namn på.  
Nytt  
Ange det nya namnet för det valda textblocket här.  
Förkortning  
I det här fältet kan Du ange en förkortning för det aktuella textblocket.  
Redigera post i litteraturförteckning  
Här redigerar du en post som har infogats i litteraturförteckningen.  
Post  
Kort beteckning  
Här ser du den korta beteckningen.  
Författare, Titel  
Här ser du postens författare och titel.  
Ändra  
Klicka här för att ändra hänvisningen till texten.  
Om du har definierat en ny datapost med kommandoknappen Ny måste du i varje fall infoga den även som post eftersom dataposten går förlorad när du stänger dokumentet annars.  
Stäng  
Stänger dialogrutan.  
Ny  
Öppnar dialogrutan Definiera litteraturpost med en tom inmatningsmask.  
Redigera  
Öppnar dialogrutan Definiera litteraturpost och visar den aktuella dataposten för redigering.  
Information om att arbeta med litteraturförteckningsposter.  
Redigera fältkommando  
Med den här funktionen öppnar du en dialogruta där du kan redigera parametrar för fältkommandon.  
I dialogrutan kan du granska och ändra det valda fältkommandot.  
Här kan du också hoppa till föregående eller nästa fältkommando i dokumentet med hjälp av två kommandoknappar och växla mellan fältkommandona av en viss typ.  
Du hittar fältkommandona lättare om du aktiverar menykommandot Visa - Fältkommandon.  
Nu visas fältnamnen och inte fältinnehållen.  
Du kan bara välja menykommandot Fältkommando... på menyn Redigera om markören står omedelbart framför ett fältkommando.  
Du kan också öppna dialogrutan för redigering av ett fältkommando genom att dubbelklicka på fältkommandot.  
Utseendet på dialogrutan avgörs av den fälttyp som är vald för tillfället, och motsvarar allmänt sett motsvarande flik i dialogrutan Fältkommandon, som Du använder för att infoga fältkommandot i fråga.  
Om Du vill redigera en DDE -länk väljer Du menykommandot Redigera - Fältkommando..., varvid dialogrutan Redigera länkar öppnas.  
Då visas dialogrutan Användardata, där Du kan göra de ändringar Du vill.  
Fälttyp  
Här ser Du det aktuella fältkommandots typ.  
Följande dialogrutselement visas bara om Du har valt tillhörande fältkommando.  
Dialogrutselement som Du inte kan aktivera, är inte tillgängliga för redigering av det aktuella fältkommandot.  
Urval  
Här visas namnet på det fält som hör till den valda fälttypen, och om flera poster föreligger kan Du välja ett annat fältkommando.  
Format  
Här kan Du ändra det aktuella fältkommandots format.  
Antalet visade alternativ bestäms av fältkommandots typ.  
När det gäller egendefinierade fält och datum - och klockslagsfält kan Du ange önskat format i dialogrutan Talformat under posten "Ytterligare format... "..  
Korrigering  
Här visas ett inställt korrigeringsvärde för sidnumret.  
Det kan Du ändra efter behov.  
Nivå  
För ett fältkommando av typ Kapitel visas här det definierade värdet på kapitelnivån, vilket Du kan ändra.  
Namn  
Här visas namnet på en fältvariabel.  
Värde  
Här står fältvariabelns aktuella värde.  
Ange ett nytt värde eller använd det förinställda.  
Villkor  
För fält som är kopplade till ett villkor visas villkoret här.  
Du kan ändra villkoret här.  
Så, annars  
För fält som är kopplade till ett villkor kan du här ändra fältinnehåll som är beroende av det villkoret.  
Hänvisning  
Här kan Du skriva eller ändra hänvisningstexten för fälttypen i fråga.  
Makronamn  
För fält som är kopplade till ett makro visas makronamnet här.  
Platshållare  
För ett fält av typen Platshållare visas platshållaren här.  
Den kan Du ändra efter behov.  
Infoga text  
Här visas den text som är kopplad till ett villkor.  
Du kan ändra en befintlig post om Du vill.  
Formel  
Om det gäller ett formelfält kan Du redigera formeln här.  
Databasurval  
Här väljer Du någon av de anmälda databaserna, om Du vill byta databas för det infogade fältkommandot.  
Du kan också välja en ny tabell eller sökning inom samma databas, som fältkommandot i fråga ska hänvisa till.  
Datapostnummer  
För ett databasfält av typen Slumpvis datapost kan Du här ändra det datapostnummer som ska infogas som fältinnehåll, om kriteriet under Villkor är uppfyllt.  
Vänsterpil  
Om Du klickar på den här kommandoknappen flyttas markören till föregående fältkommando av samma typ.  
Knappen är tillgänglig bara om det finns flera fältkommandon av samma typ i dokumentet.  
Föregående fältkommando  
Högerpil  
Om Du klickar på den här kommandoknappen flyttas markören till nästa fältkommando av samma typ.  
Knappen är tillgänglig bara om det finns flera fältkommandon av samma typ i dokumentet.  
Nästa fältkommando  
Redigera fotnot  
Med det här kommandot kan du redigera den aktuella fotnoten.  
Dialogrutan Redigera fotnot ger samma möjligheter som dialogrutan Infoga fotnot.  
Här kan du ändra alla inställningar som du gjorde när du infogade fotnoten.  
Du kan använda kommandot Fotnot... på menyn Redigera bara om textmarkören står omedelbart framför eller på fotnotstecknet.  
Du ändrar texten i fotnoten helt enkelt genom att först klicka i fotnotstexten nederst på sidan (eller sist i dokumentet) och sedan redigera texten.  
Du kan hoppa från fotnotsankaret till fotnoten med musen.  
Den blir då till en hand med utsträckt pekfinger.  
Om Du klickar nu, hoppar markören till själva fotnotstexten.  
Du kommer tillbaka till fotnotsankaret med tangenten PageUp (PgUp).  
Numrering  
Här väljer Du typ av fotnotsnumrering för den aktuella fotnoten.  
Automatisk  
Tecken  
...  
Det är lätt att ändra ett fotnotsteckens formatering och teckensnitt.  
Du kan också använda motsvarande formateringsfunktioner på objektlisten.  
Typ  
Här väljer Du om det gäller en fotnot eller slutnot.  
Fotnot  
Med det här alternativet kan Du växla från slutnoter till fotnoter.  
Slutnot  
Med det här alternativet kan Du växla från fotnoter till slutnoter.  
Vänsterpil  
Om Du klickar på den här kommandoknappen placeras markören i föregående fotnot.  
Föregående fotnot  
Högerpil  
Om Du klickar på den här kommandoknappen placeras markören i nästa fotnot.  
Nästa fotnot  
Redigera förteckningspost  
Här kan Du redigera förteckningsposter.  
Den här funktionen kan Du bara använda om markören står i eller omedelbart framför en förteckningspost.  
De förteckningsposter som har infogats i texten med Infoga - Förteckningar - Post... redigeras.  
Markering  
I det här området redigerar Du förteckningsposten.  
Förteckning  
I det här fältet visas den aktuella postens förteckningstyp.  
Du kan inte ändra en posts typ.  
Om Du trots det vill göra det, måste Du först radera posten och lägga in den under en ny typ.  
Post  
De tillägg som Du gör här visas bara i förteckningen, inte i löptexten.  
Här kan Du t ex utvidga en sakordsförteckningspost med kommentarer, t ex "Övrigt, se även Allmänt".  
Sorteringskod 1  
Om Du vill skapa ett register där sakorden är uppställda på flera nivåer anger Du här "övertermen" på den högsta nivån, eller också väljer Du den "överterm "som det aktuella sakordet ska underordnas.  
Sorteringskod 2  
Om Du vill skapa ett register där sakorden är uppställda på flera nivåer, anger Du här "övertermen" på nivå två, eller också väljer Du den "överterm "som det aktuella sakordet ska underordnas.  
Nivå  
Om Du vill dra in de poster i innehållsförteckningens som motsvarar kapitelnivå åt höger, anger Du önskad nivå här.  
Radera  
Med den här kommandoknappen tar Du bort den aktuella förteckningsposten.  
Det är bara posten i förteckningen som försvinner, inte motsvarande markerade ord i löptexten.  
De efterstående riktningspilarna visas bara om det finns flera identiska förteckningsposter i dokumentet.  
Stoppil åt vänster  
Leder till föregående förteckningspost av samma typ och med samma innehåll i dokumentet.  
Stoppil åt vänster  
Stoppil åt höger  
Leder till nästa förteckningspost av samma typ och med samma innehåll i dokumentet.  
Stoppil åt höger  
De efterstående riktningspilarna visas bara om det finns flera identiska förteckningsposter i dokumentet.  
Vänsterpil  
Leder till föregående förteckningspost av samma typ i dokumentet.  
Vänsterpil  
Högerpil  
Leder till nästa förteckningspost av samma typ i dokumentet.  
Högerpil  
Du kan också snabbt hoppa till olika förteckningsposter i dokumentet med hjälp av navigationslisten.  
Redigera områden  
Här kan du redigera egenskaperna för områdena som är definierade i dokumentet.  
Du kan bara använda kommandot om du dessförinnan har infogat minst ett område.  
Dialogrutan Redigera områden är uppbyggd som fliken Område i dialogrutan Infoga område, som Du öppnar med menykommandot Infoga - OmrÃ¥de...  
Dessutom hittar Du följande alternativ i Redigera områden.  
Område  
I listrutan Område markerar du namnet på det område som ska redigeras eller namnen i en multimarkering, eller också skriver du områdesnamnet i textfältet Område.  
På statuslisten nere till höger kan du se i vilket område textmarkören för tillfället står.  
Till vänster intill områdesnamnet anges med små symboler om området är skyddat (ett stängt hänglås), oskyddat (öppet hänglås) eller om det är synligt, alltså inte dolt (små glasögon).  
De här egenskaperna kan Du ställa in för flera områden samtidigt.  
Alternativ  
Med den här kommandoknappen öppnar du dialogrutan Alternativ där du kan redigera kolumner, bakgrund, fot - och slutnoter.  
Om området är skyddat med ett lösenord måste du ange lösenordet först.  
Upphäv  
Texten i det markerade området blir en normal text.  
Linjal  
Med det här kommandot kan du visa respektive dölja linjaler.  
Om menykommandot är markerat, visas linjalerna till vänster och ovanför arbetsområdet.  
Som förinställning visar %PRODUCTNAME Writer bara den horisontella linjalen ovanför arbetsområdet.  
Om du vill att även den vertikala linjalen ska visas, väljer du Verktyg - Alternativ - Textdokument - Vy och markerar rutan för den vertikala linjalen.  
Linjalerna visar indelningen av arbetsområdet i det aktuella dokumentet.  
På den horisontella linjalen visas dessutom tabbstoppen.  
Arbetsområdet anges på linjalen av det ljusa området.  
Om Du vill ändra indraget från vänster på den horisontella linjalen kan Du göra det med markeringen till vänster på linjalen.  
Om Du vill flytta högermarginalen, gör Du det med markeringen till höger på linjalen.  
Om Du vill infoga ett tabbstopp i dokumentet klickar Du på linjallisten.  
Den tabbtyp som visas intill linjalen infogas där Du klickar.  
Genom att klicka på symbolen till vänster om linjalen växlar Du mellan de olika tabbtyperna.  
Med den övre trekanten på linjallisten kan Du göra ett indrag av första raden i ett enskilt stycke respektive kontrollera avståndet från marginalen för rader som redan är indragna.  
Den undre trekanten till höger anger dokumentets högermarginal.  
Om Du vill ändra högermarginalen, placerar Du trekanten där Du vill att den nya marginalen ska vara.  
Om dokumentet innehåller en tabell och markören står i denna, visas kolumnbredderna med skiljelinjer på linjalen.  
Den aktuella kolumnen markeras på linjalen med vänster och höger begränsningstecken.  
På så vis kan Du ange indrag till vänster och höger för kolumnen.  
Dessutom kan Du ändra kolumnbredden med hjälp av linjalen.  
Ställ muspekaren på linjallisten på den kolumnbredd som är markerad med en skiljelinje.  
Muspekaren förvandlas till en dubbelpil.  
Klicka på skiljelinjen, håll musknappen nedtryckt och dra linjen till önskad position.  
Kolumnbredden ställs direkt in på den nya bredden.  
Om Du vill att kolumnbredderna ska bibehålla sina inbördes proportioner när Du ändrar en kolumn, håller Du ned Kommando Ctrl -tangenten när Du ändrar.  
Alla kolumner efter den kolumn som ändras förskjuts i förhållande till sina bredder.  
Om grafiska objekt, ramar eller andra objekt är aktiva i dokumentet, visas respektive storlek på linjalerna.  
För sidhuvud och sidfötter bibehåller den horisontella linjalen sin disposition, medan den vertikala linjalen visar radhöjden.  
Om du vill ändra en tabulator, placerar du muspekaren på den och öppnar snabbmenyn.  
Alternativt kan du dubbelklicka på tabulatorn.  
Dialogrutan motsvarar den som öppnas om du väljer menykommandot Format - Stycke - Tabulator visas.  
Om du dubbelklickar på linjallisten öppnas en dialogruta som motsvarar menykommandot Format - Stycke.  
Måttenheten för linjalerna väljer du i dialogrutan Verktyg - Alternativ - Textdokument - Vy.  
Där ställer du också in avståndet för tabbar, som annars är förinställda på mått som gäller tills du ersätter dem med egna tabbar.  
Du kan också ställa in tabbar, indrag, marginaler, kolumner och mått på markerade objekt med musen och ställa in linjalernas måttenheter via snabbmenyn.  
Om du vill radera en tabulator klickar du på den och drar den med nedtryckt musknapp nedåt från linjallisten.  
Textbegränsningar  
Med det här kommandot kan du visa eller dölja textbegränsningar.  
Textbegränsningar är linjer och som visar marginaler, ramar, objektkanter o.s.v. på bildskärmen, men som inte skrivs ut.  
Om menykommandot är markerat är visningen av textbegränsningar aktiverad.  
Huruvida textbegränsningarna visas eller inte har ingen betydelse för det utskrivna dokumentets utseende.  
De är bara till för att underlätta överblicken över dokumentet på bildskärmen.  
Markeringar  
Med det här kommandot sätter du på eller stänger av visningen av markeringar i texten.  
Exempel på sådana markeringar är fasta mellanrum, användardefinierade bindestreck, förteckningsposter, fotnotstecken och fält.  
Följande textelement berörs av markeringar:  
Element  
Visning  
Fast mellanrum  
Fast mellanrum, som alltid håller ihop ord, har grå bakgrund.  
Användardefinierade bindestreck  
Användardefinierade bindestreck visas i texten.  
Förteckningsposter  
Förteckningsposter visas med grå bakgrund.  
Bakgrundsfärg för fotnoter  
Fotnotsnummer visas med grå bakgrund.  
Bakgrundsfärg för fält  
Infogade fält visas med grå bakgrund.  
När du ska definiera vilka av ovannämnda textelement som ska visas väljer du Verktyg - Alternativ - Textdokument - Formateringshjälp.  
Förutom markeringarna kan du även låta kontrolltecknen visas.  
Du använder ikonen Kontrolltecken på / av på verktygslisten.  
Fältkommandon  
Här växlar du mellan visning av namn på fältkommandon och deras innehåll.  
I annat fall visas själva innehållet i fältkommandona.  
Fältkommandonas namn visas alltid, däremot visas i många fall inte deras innehåll.  
Mer information om fältkommandon finns under Infoga - Fältkommando.  
Den här funktionen kan du även aktivera och inaktivera i den dialogruta som du öppnar med Verktyg - Alternativ... - Textdokument - Vy under "Visa - Fältnamn".  
Om du skriver ut ett dokument när visningen av fältkommandon som fältnamn är aktiverad visas först en dialogruta.  
Här kan du välja om du vill skriva ut dokumentet med fältnamn (Ja), om du vill skriva ut det utan fältnamn, alltså med värdena respektive innehållet i fältkommandona (Nej), eller om du vill avbryta åtgärden.  
Kontrolltecken  
Välj den här funktionen när du vill sätta på eller stänga av visningen av kontrolltecken i texten.  
Några exempel på kontrolltecken är radbrytning, tabulatorer och blanksteg.  
Kontrolltecknen visar styckeslut, tabbar och blanksteg.  
Styckeslut utgörs av ett synlig stycketecken, tabbar visas med en liten högerpil, och ett blanksteg med en punkt.  
Om det finns en bock framför menyalternativet, visas kontrolltecknen som finns i dokumentet i arbetsområdet.  
Detta är till hjälp om du t.ex. vill kopiera delar som börjar eller slutar med sådana tecken och klistra in dem på en annan plats.  
Särskilt viktiga är stycketecknen, eftersom de innehåller formateringsinformationen om det följande stycket.  
Om du raderar ett stycketecken, får följande stycke samma formatering som det föregående.  
Om du raderar stycketecknet omedelbart framför en tabell, raderas hela tabellen.  
När du ska definiera vilka kontrolltecken som ska visas, väljer du Verktyg - Alternativ - Textdokument - Formateringshjälp.  
Visningen av kontrolltecken på bildskärmen påverkar inte utskriften.  
Onlinelayout  
Med kommandot Onlinelayout ser du %PRODUCTNAME Writer-dokumentet som om det rörde sig om ett HTML-dokument.  
Den här funktionen är särskilt praktisk när du skapar dokument för Internet.  
I onlinelayouten visas dokumentet med dokumentmallen html.stw.  
I den här vyn kan Du använda en mycket lång sida, så att den som tittar på den som Internetsida endast i sällsynta fall behöver störas av sidbrytningar.  
Om Du tidigare har öppnat flera visningar (på menyn Fönster - Nytt fönster), stängs övriga fönster när Du går över till onlinelayout.  
Utskriftslayout  
Använd det här kommandot om du vill se hur layouten ser ut när dokumentet är utskrivet.  
Kommandot Visa - Utskriftslayout är bara tillgängligt när ett HTML-dokument är öppet.  
Dolda stycken  
Med det här kommandot sätter du på och stänger av visningen av dolda stycken på skärmen.  
Du kan även aktivera den här funktionen via rutan Dolda stycken under Verktyg - Alternativ - Textdokument - Formateringshjälp.  
Dolda stycken är stycken vars visning du gör beroende av ett villkor med hjälp av fältkommandot "Dolt stycke".  
Om villkoret uppfylls, döljs stycket och finns inte med på utskriften.  
Ifall villkoret inte uppfylls, döljs stycket inte och skrivs alltså ut.  
I det här fallet spelar det ingen roll om alternativet för visning av dolda stycken har markerats eller inte, eftersom den här kryssrutan bara styr visningen på bildskärmen.  
När ett dolda stycken döljs så döljs även deras fotnoter och ramar som är bundna till tecken.  
Infoga brytning  
Med den här funktionen infogar du en manuell rad-, kolumn - eller sidbrytning vid markörens position.  
Typ  
Här väljer Du typ av brytning.  
Radbrytning  
Den text som står till höger om markören flyttas till början av nästa rad, men något nytt stycke påbörjas inte.  
Du åstadkommer samma sak genom att trycka på Skift+Retur.  
Kolumnbrytning  
Texten till höger om markören flyttas till början av nästa kolumn.  
En sådan kolumnbrytning markeras genom att den nya kolumnen får en blå överkant.  
Sidbrytning  
Texten till höger om markören flyttas till början av nästa sida.  
En sådan sidbrytning markeras genom att den nya sidan får en blå överkant.  
Du kan infoga en sidbrytning genom att trycka på Kommando Ctrl +Retur.  
Om Du vill kunna använda en annan sidformatmall på nästa och följande sidor måste Du dock infoga den manuella sidbrytningen med menykommando, inte med kortkommando.  
Formatmall  
Vid en sidbrytning kan Du här ange sidformatmall för nästa sida.  
Ändra sidnummer  
Om den automatiska sidnumreringen på sidan efter sidbrytningen ska ändras, markerar Du den här kryssrutan.  
Ange sidnumret i fråga i det nedre rotationsfältet.  
Sidnummer  
Här anger Du det nya sidnummer som ska gälla efter den manuella brytningen.  
Med menykommandot Visa - Styrtecken visar Du de manuellt infogade radbrytningarna.  
> Infoga omrÃ¥de  
Med den här funktionen infogar du ett område vid markörens position.  
Området kan behandlas separat från normaltexten och på det här sättet kan du dölja textavsnitt, arbeta med olika kolumnindelningar per sida eller skydda stycken mot ändringar.  
Dessutom kan du koppla visningen av ett område till vissa villkor.  
Vidare kan du skapa en länk för ett område till en annan fil eller ett namngivet område i den andra filen eller skapa den via DDE.  
Om du ska redigera infogade områden väljer du menykommandot Format - Områden....  
%PRODUCTNAME skapar området för markerade textställen.  
Om ingen text är markerad, infogas en styckebrytning och definieras som område.  
Följande flikar visas:  
Infoga  
Med den här kommandoknappen infogar du området med de inställningar som du har gjort på den plats i dokumentet där markören står.  
Område  
Här ger du området ett namn och ställer in alternativen.  
Nytt område  
Det börjar alltid med Område1.  
Länk  
Länka  
Om du markerar den här rutan, kan du länka ett område i ditt dokument till ett annat område i en annan fil.  
DDE  
Om du har aktiverat rutan Länka, kan du också skapa en länk via DDE.  
I så fall markerar du rutan DDE och skriver in önskat DDE-kommando i textfältet DDE-kommando.  
Syntaxen för ett DDE-kommando ser i allmänhet ut så här: "<Server> <Topic> <Item>".  
Server är DDE-namnet på det program som tillhandahåller data.  
Topic är den plats, där Item är placerat, dvs för det mesta filnamnet, och Item är det enskilda objekt som tillhandahålls.  
Två exempel:  
Du vill infoga området med namnet Område1 från %PRODUCTNAME -textdokumentet abc.sdw via DDE.  
DDE-kommandot lyder: "soffice x:\abc.sdw Område1".  
Du vill infoga den första cellens innehåll från en MS-Excel-tabell i filen abc.xls.  
DDE-kommandot lyder: "excel x:\[abc.xls]Tabell1 z1s1".  
Om Du kopierar motsvarande element och sedan infogar urklippets innehåll som DDE-länk med kommandot Redigera - Klistra in innehåll..., visas syntaxen om Du väljer menykommandot Redigera - Fältkommando....  
Filnamn / DDE-kommando  
Skriv in filens sökväg och namn här eller, om DDE är markerat, DDE-kommandot.  
...  
Med hjälp av den här kommandoknappen hittar du en fil.  
Den aktiveras bara om rutan Länka är markerat.  
Område  
Här kan Du markera ett område för länkning i den angivna filen.  
Genom länkningen visas innehållet i den länkade filen, eller det markerade området i filen, i det aktuella dokumentets markerade område.  
När dokumentet laddas på nytt tillfrågas Du om länkarna ska uppdateras.  
Skrivskydd  
Skyddat / Skydda  
Om innehållet i området inte ska ändras eller redigeras mer, markerar du den här rutan.  
På så vis förhindrar du t.ex. att element i området redigeras eller flyttas av misstag.  
Med lösenord  
I kombination med ett lösenord kan du också förhindra att området ändras av obehöriga personer.  
...  
Klicka här om du vill ange ett lösenord.  
Dölj  
Dölj  
Om det markerade området inte ska visas, markerar du den här rutan.  
På det här sättet kan du t.ex. temporärt förhindra att delar av dokumentet visas eller skrivs ut eftersom du inte vill att de ska vara läsbara ännu, men som du ändå vill ta med i dokumentet av organisatoriska skäl.  
Innehållet i dolda områden (t.ex. grafik) visas i grått i Navigator.  
Tipshjälpen visar texten "dolt".  
Du kan upphäva de dolda områdena under Format - Områden  
Med villkor  
Om du vill att området bara ska visas eller skrivas ut när vissa villkor uppfylls, klickar du i det här textfältet och anger villkoret för visningen av området.  
Det går bara att ändra ett villkor om rutan Dölj är markerad.  
Villkor  
Ange här det villkor som ska uppfyllas för att området ska döljas.  
Om villkoret är sant (TRUE), döljs området, och om det är falskt (FALSE), döljs det inte.  
Villkoren är logiska uttryck, som t.ex. "TILLTAL EQ Mr. ".  
Här kan du t.ex. ange att i ett standardbrev (kopplad utskrift) ska ett område, vars tillhörande databas innehåller fältet "Tilltal "med innehållet "Mr .", "Ms." eller "Sir or Madam", bara visas eller skrivas ut om tilltalet är lika med "Mr. ".  
Eller så definierar du en fältvariabel x och sätter dess värde till 1.  
Ange sedan följande villkor för Dölj: "x eq 1" i det här fältet.  
Det definierade området visas inte förrän du tilldelar fältvariabeln x ett annat värde.  
Mer information om fältkommandon och syntaxen för villkor hittar du på respektive ställe i hjälpen.  
Infoga fotnot  
Med den här funktionen infogar du en fotnot.  
Du kan välja mellan automatisk numrering och en fotnotsvisning som du kan definiera själv, och du kan bestämma om det ska vara en fotnot eller en slutnot.  
Följande beskrivning av fotnoter gäller även för slutnoter.  
Slutnoter är fotnoter som samlas vid dokumentets slut i stället för längst ner på sidan.  
Numrering  
Här väljer du typ av fotnotsnumrering för fotnoten som ska infogas.  
Automatisk  
Aktivera det här alternativfältet om du vill använda den automatiska fotnotsnumreringen.  
Då används inställningarna som du har gjort under Verktyg - Fotnoter... i dialogrutan Fotnotsinställning.  
Tecken  
Med det här alternativet kan du för den aktuella fotnoten ange ett tecken som du skriver i textfältet intill.  
Det kan vara en bokstav eller ett nummer.  
Du kan också använda ett specialtecken med kommandoknappen nedanför.  
...  
Om Du klickar på den knappen öppnas en dialogruta där Du kan välja ett specialtecken.  
Om Du gör det, visas tecknet i textfältet.  
Typ  
Här väljer du om du ska infoga en fotnot eller en slutnot.  
Medan du för fotnoter kan välja om de ska infogas nedtill på sidan eller i slutet av dokumentet, samlas slutnoter alltid i slutet av dokumentet.  
Slutnoter och fotnoter numreras separat från varandra.  
Fotnot  
Välj det här alternativet om du vill infoga en fotnot.  
Slutnot  
Välj det här alternativet om du vill infoga en slutnot.  
Information om att arbeta med fotnoter.  
Infoga bokmärke  
Med den här funktionen infogar du ett bokmärke där markören står.  
Bokmärken listas med sina namn i Navigator, och därifrån kan du direkt hoppa till dem.  
I HTML-dokument ser bokmärken ut som ankare som du kan hoppa till med hjälp av hyperlänkar.  
Du kan använda bokmärken till att hoppa till bestämda platser i texten med Navigator.  
Om texten innehåller bokmärken, indikeras detta i Navigator med små plustecken bredvid de poster där bokmärkena finns.  
Om Du klickar med musen på ett plustecken eller dubbelklickar på en bokmärkespost i Navigator, öppnas en lista över bokmärkena.  
Om Du dubbelklickar på en bokmärkespost i Navigator, flyttas markören i dokumentet till bokmärkets plats.  
Du kan också öppna den här popup-menyn genom att klicka med höger musknapp i fältet Sidnummer på statuslisten.  
Om Du sedan klickar en gång på bokmärkets namn, flyttas textmarkören till önskad plats.  
Bokmärken  
I det övre textfältet anger Du det nya bokmärkets namn.  
I den undre listrutan listas de bokmärken som finns i dokumentet.  
Om Du klickar på ett bokmärke på listan förs motsvarande namn in i textfältet, där Du kan redigera det.  
Dock får Du inte använda följande tecken: /\ @: *? ";,. #  
Radera  
Om Du vill ta bort ett bokmärke, markerar Du det i listrutan i dialogrutan Infoga bokmärke och klickar sedan på Radera.  
Då raderas bokmärket utan att Du ombeds bekräfta det.  
Bildtext  
Med den här funktionen infogar du bildtexter och automatiska numreringar.  
Det kan vara bildtexter till tabeller, ramar, grafikobjekt, textramar eller ritobjekt.  
Kommandot finns också i respektive snabbmeny.  
Egenskaper  
Ovanför fälten där du gör dina inställningar visas den aktuella numreringen av bildtexten bredvid den aktuella kategorin.  
Kategori  
Här visas vilken styckeformatmall som gäller för det markerade objektet.  
Varje objekttyp har som standard en egen styckeformatmall.  
Illustration, Tabell, Text och Teckning.  
Du kan naturligtvis definiera en egen styckeformatmall eller använda en annan mall för bildtexterna till dina objekt.  
Det gör du helt enkelt genom att ange den önskade styckeformatmallen i fältet Kategori.  
Den text som du anger under Kategori förs över till bildtexten.  
Om du t.ex. vill använda texten "Fig 1" som bildtext i stället för "Figur 1", skriver du helt enkelt "Fig "i stället för "Figur".  
En kopia av mallen skapas då med det här nya namnet.  
Numrering  
Välj numreringstyp här.  
Bildtext  
Här skriver du bildtexten.  
Den inskrivna texten visas direkt efter numreringen.  
Om du t.ex. vill att dina objekt ska beskrivas enligt mönstret "Objekt 1:  
Text ", skriver du under Bildtext först ett kolon, sedan ett blanksteg och slutligen den text som ska höra till objektet.  
Position  
Här kan du i förekommande fall ange hur bildtexten ska placeras.  
Objekttypen avgör om den här funktionen är tillgänglig och vilka alternativ som i så fall finns.  
Överta inramning och skugga  
Om du markerar den här rutan utvidgas inramningen och skuggningen till bildtextområdet.  
Objektnamn  
Här ger du objektet det namn som det ska ha i t.ex. Navigator.  
Alternativ  
Sekvensalternativ  
Här ställer du in den nivå, där nummersekvensen (t.ex. i en bildtext) ska börja om på 1 när nivån ändras.  
Numrering kapitelvis  
I det här området anger du hur numreringen av kapitel ska börja om.  
Nivå  
Här väljer du den rubrik - respektive kapitelnivå vid vilken numreringen ska börja om när nivån ändras i dokumentet.  
Skiljetecken  
Ange här det tecken som ska stå mellan numret på överskrifts - respektive kapitelnivån och numret på det rubrikförsedda objektet.  
Kuvert  
Med den här funktionen skapar du ett kuvert.  
Du definierar kuvertstorlek, justering av kuvertet vid utskrift och avsändar - och mottagaradress.  
Nytt dok.  
Om du klickar på den här kommandoknappen skapas ett nytt dokument enligt uppgifterna som du har angett i dialogrutan.  
Infoga  
Klicka på den här kommandoknappen när Du inte vill skriva ut det definierade textområdet på ett kuvert utan i stället infoga det i dokumentet.  
Då infogas en extrasida framför den aktuella sidan som har sidformatmallen "Kuvert".  
Kuvert  
Här anger du data för mottagare och avsändare på kuvertet.  
Du kan hämta motsvarande fält i en datakälla.  
Mottagare  
Här anger du mottagaren.  
Du kan välja mellan att skriva texten direkt resp. att kopiera den från urklippet, eller att placera markören där texten ska stå och sedan välja ett datafält från en datakälla vars innehåll ska klistras in där markören står.  
Texformateringar, t.ex. fetstil, kan du göra efteråt i texten på kuvertsidan.  
Avsändare  
Markera den här rutan om kuvertet ska ha ett område för avsändaren.  
Ange en avsändare i textfältet.  
Avsändardata hämtas från användardata, men du kan ändra dem.  
Databas  
I det här kombinationsfältet väljer du den databas som innehåller uppgifterna om mottagaren.  
Tabell  
Här väljer du den databastabell där du vill hämta underlag för mottagaruppgifterna.  
Databasfält  
Välj ett databasfält i det kombinationsfält som hör till den utvalda databasen.  
Om du klickar på pilen, infogas databasfältets innehåll i fältet Mottagare där markören står.  
Format  
Här väljer du placering och format för avsändar - och mottagarfält.  
Även formatet på kuvertet som ska skrivas ut ställer du in här.  
Mottagare  
Här väljer du placeringen och formatet för mottagarfältet på kuvertet.  
Placering  
I det här området bestämmer du samtliga egenskaper för placeringen av mottagarområdet på kuvertet.  
från vänster  
I det här rotationsfältet ställer du in var mottagarområdet ska börja i förhållande till kuvertets vänsterkant.  
uppifrån  
I det här rotationsfältet ställer du in var mottagarområdet ska börja i förhållande till kuvertets överkant.  
Format Redigera  
Den här popupmenyn öppnar Du när Du ska byta mellan redigering av tecken - och styckeegenskaper för styckeformatmallen "Mottagare".  
Tecken...  
När du väljer det här kommandot på undermenyn visas en dialogruta med följande flikar:  
Teckensnitt, Teckeneffekt, Hyperlänk, Bakgrund, Position och om stödet för asiatiska språk är aktiverat Asiatisk layout  
Under de här flikarna väljer du teckenformatering för texten i kuvertets mottagarfält.  
Stycke...  
När du väljer det här kommandot på undermenyn visas en dialogruta med följande flikar:  
Indrag och avstånd, Justering, Textflöde, Tabulator, Anfanger, Inramning, Bakgrund och om stödet för asiatiska språk är aktiverat Asiatisk typografi.  
Under de här flikerna väljer du styckeformatering för texten i kuvertets mottagarfält.  
Avsändare  
Här väljer du placeringen och formatet för avsändarfältet på kuvertet.  
Placering  
I det här området bestämmer du alla egenskaper för placeringen av avsändarområdet på kuvertet.  
från vänster  
I det här rotationsfältet ställer du in var avsändarområdet ska börja i förhållande till kuvertets vänsterkant.  
uppifrån  
I det här rotationsfältet ställer du in var avsändarområdet ska börja i förhållande till kuvertets överkant.  
Format Redigera  
Den här popupmenyn öppnar Du när Du ska byta mellan redigering av tecken - och styckeegenskaper för styckeformatmallen "Avsändare".  
Tecken...  
När du väljer det här kommandot på undermenyn visas en dialogruta med följande flikar:  
Teckensnitt, Teckeneffekt, Hyperlänk, Bakgrund, Position och om stödet för asiatiska språk är aktiverat Asiatisk layout.  
Där väljer Du teckenformatering för texten i kuvertets avsändarfält.  
Stycke...  
När Du väljer det här undermenyalternativet visas en dialogruta med följande flikar:  
Indrag och avstånd, Justering, Textflöde, Tabulator, Anfanger, Inramning, Bakgrund och om stödet för asiatiska språk är aktiverat Asiatisk typografi.  
Där väljer Du styckeformatering för texten i kuvertets avsändarfält.  
Storlek  
Här väljer Du kuvertets format.  
Du väljer antingen något av de förinställda formaten eller så anger Du värdena för bredd och höjd.  
Format  
I den här listrutan väljer Du kuvertformat bland ett antal förinställda standardiserade kuvertformat.  
Fälten Bredd och Höjd får motsvarande värden.  
Dessa värden kan Du alltid ändra.  
Bredd  
Här ställer Du in kuvertets bredd.  
Höjd  
Här ställer Du in kuvertets höjd.  
Skrivare  
Här anpassar du utskriftsposition och -justering till skrivaren som du använder.  
Se efter i skrivarens dokumentation hur Du måste lägga in kuverten för att de ska matas igenom skrivaren på rätt sätt.  
Beroende på skrivarmodell kan det hända att kuverten måste läggas an mot vänster sida, mot höger sida eller placeras i mitten; och i vissa skrivare måste de placeras med utskriftssidan nedåt, i andra med den uppåt.  
Liggande till vänster  
Kuvertet läggs in mot fackets vänstra sida och blir liggande.  
Liggande i mitten  
Kuvertet läggs in i mitten av facket i liggande riktning.  
Liggande till höger  
Kuvertet läggs in mot fackets högra sida i liggande riktning.  
Stående till vänster  
Kuvertet läggs in mot fackets vänstra sida i stående riktning.  
Stående i mitten  
Kuvertet läggs in i mitten av facket i stående riktning.  
Stående till höger  
Kuvertet läggs in mot fackets högra sida i stående riktning.  
Skriv ut uppifrån  
Kuvertet läggs in med den sida uppåt där texten ska hamna.  
Skriv ut nedifrån  
Kuvertet läggs in med den sida nedåt där texten ska hamna.  
Åt höger  
Här fininställer Du den horisontella positionen för det område som ska skrivas ut.  
Nedåt  
Här fininställer Du den vertikala positionen för det område som ska skrivas ut.  
Aktuell skrivare  
Här visas namnet på den aktuella skrivaren.  
Du växlar aktuell skrivare i operativsystemet.  
Ställ in...  
Den här kommandoknappen öppnar dialogrutan Skrivarinställning.  
Här kan Du, beroende på vilken skrivare Du använder, göra fler inställningar, t ex för använt pappersformat och orientering.  
Fältkommandon  
Den här funktionen öppnar en dialogruta med vars hjälp du infogar ett fältkommando.  
I dialogrutan kan du välja alla tillgängliga fältkommandon.  
Infoga  
Om Du klickar på den här kommandoknappen infogar Du det markerade fältkommandot där markören står i dokumentet.  
Dialogrutan är fortfarande öppen.  
Om Du vill infoga ytterligare ett fältkommando, behöver Du bara sätta markören i önskad position i dokumentet och sedan välja nästa fältkommando i dialogrutan.  
Dokument  
Dokumentfält används till att infoga innehåll som har en direkt relation till det aktuella dokumentet.  
Utöver dokumentets specifika kännetecken, t.ex. filnamn, dokumentmall och statistiska uppgifter, kan dokumentfält även innehålla användardata, datum och klockslag.  
När datum - och tidsfält importeras och exporteras i HTML-format, gäller speciella %PRODUCTNAME -format.  
Fälttyp  
Här väljer du fälttyp.  
Du kan välja bland följande fälttyper:  
Fälttyp  
Betydelse  
Avsändare  
Infogar fält med uppgifter om användaren.  
Fältinnehållet registrerades vid installationen, men du kan ändra det i efterhand under Verktyg - Alternativ - %PRODUCTNAME - Användardata.  
Användare  
Infogar användarnamn eller initialer.  
Du kan ändra uppgifterna under Verktyg - Alternativ - %PRODUCTNAME - Användardata.  
Filnamn  
Infogar filnamn och / eller sökväg för det aktuella dokumentet och filnamnet utan filnamnstillägg.  
Datum  
Infogar aktuellt datum.  
Datumet kan antingen inte ändras längre (datum fast) eller uppdateras automatiskt (datum var.).  
Du väljer datumformat under Format.  
Dokumentmall  
Infogar filnamnet och / eller katalogsökvägen för den aktuella dokumentmallen samt filnamnet utan filnamnstillägg.  
De använder namnen som visas för mallförvaltning i %PRODUCTNAME i dialogrutan Dokumentmallar.  
Kapitel  
Infogar kapitelnummer och / eller kapitelnamn.  
Sida  
Infogar sidnumret för den aktuella, föregående eller följande sidan.  
Statistik  
Infogar statistiska uppgifter om dokumentets innehåll, dvs sidor, stycken, ord, tecken, tabeller, grafiska objekt och andra objekt.  
Klockslag  
Infogar aktuell systemtid.  
Klockslaget är antingen låst (klockslag fast) eller uppdateras om Du uppdaterar fältet med F9 (klockslag var.).  
Följande textfält visas bara eller kan bara aktiveras om Du har valt motsvarande fälttyp.  
Urval  
Välj ett fältkommando här.  
Det finns en beskrivning av hur du arbetar med sidformatmallar och sidnummer här.  
För fältkommandon av typen Sida har du följande alternativ att välja mellan:  
Fältkommando  
Funktion  
Föregående sida  
Infogar sidnumret för föregående sida.  
Nästa sida  
Infogar sidnumret för nästa sida.  
Sidnummer  
Infogar sidnumret för den aktuella sidan.  
Under Format kan Du välja önskat visningsformat för sidnummer.  
Om Du väljer formatet Text kan Du ange en egen text i textfältet Värde.  
Under Korrigering kan du ange en korrigeringsfaktor, t.ex. +1 eller -1, med vilken det aktuella sidnumret ändras i visningen.  
Du behöver den här funktionen om t.ex. numret på följande sida (korrigeringsvärde +1) ska stå i slutet av varje sida.  
Det beräknade sidnumret måste existera i dokumentet för att fältinnehållet ska infogas.  
Sista sidan i dokumentet visar därför automatiskt inget nummer för någon följande sida.  
Noll kan inte visas.  
Eftersom den beräknade sidan även måste finnas i dokumentet, så medför t ex korrigeringsvärdet -1 för funktionen "Föregående sida" att det är först fr o m sida 3 som resultatet blir meningsfullt.  
Använd då kommandot Infoga - Manuell brytning... och byt på så vis till en ny sidformatmall.  
Om Du håller tangenten Kommando Ctrl nedtryckt samtidigt som Du dubbelklickar på en post, så infogas denna direkt i dokumentet.  
Format  
Här väljer du formatet i vilket fältkommandot ska infogas.  
För datum - och klockslagsfält kan du, förutom de förinställda formaten, definiera ett eget format om du klickar på posten "Ytterligare format...".  
Med det här alternativet öppnar du dialogrutan Talformat.  
När Du väljer alternativet "Kapitelnummer utan skiljetecken" för ett kapitelfält, utelämnas de skiljetecken som Du har angett under Verktyg - Kapitelnumrering....  
För referensfält kan Du välja kapitelnumret som Format.  
Då visas det refererade objektets kapitelnummer i referensen.  
Om denna kapitelnivå inte är numrerad, så letar %PRODUCTNAME Writer i de överordnade nivåerna efter en nivå med numrering och infogar dess kapitelnummer.  
Om du infogar en numrering eller punktuppställning i ett stycke på en sida, d.v.s. direkt i anslutning till en text, så tilldelas numreringen eller punktuppställningen stycket.  
När du refererar till nummersekvenser kan du välja i vilket format det ska ske.  
Du kan bland annat välja följande:  
Kategori och nummer  
Formatet omfattar allting från styckets början till nummersekvensfältets slut.  
Bildtext  
Formatet omfattar texten efter nummersekvensfältet fram till stycketecknet.  
Nummer  
Detta format omfattar bara referensnumret.  
Nivå  
Här kan Du ange den önskade nivån för ett fältkommando av typen Kapitel.  
Korrigering  
Här kan du mata in det önskade korrigeringsvärdet för sidnumret för ett fältkommando som anger ett sidnummer.  
På det här sättet går det t.ex. att visa numret för den följande sidan på en sida.  
Korrigering i dagar / - minuter  
Här kan Du mata in ett önskat korrigeringsvärde för ett fältkommando som anger ett datum eller ett klockslag.  
Värde  
Här läggs fältinnehållet in vid fält som du själv definierar.  
Det här textfältet är bara tillgängligt för dokumentfält om du vill mata in numret på föregående eller nästa sida i textformat vid fältkommandon av typen sida.  
Referenser  
Här infogar du referenser resp. korshänvisningar i det aktuella dokumentet.  
Referenser är korshänvisningar inom samma dokument eller inom ett samlingsdokuments deldokument.  
Fördelen med att infoga en korshänvisning som fältkommando är att du inte måste anpassa hänvisningarna manuellt så snart du ändrar något i dokumentet.  
Du behöver bara uppdatera fältkommandona med F9, så stämmer korshänvisningarna igen.  
Fälttyp  
Betydelse  
Sätt referens  
Sätter målet för en korshänvisning.  
Under Namn anger Du en beteckning för referensen.  
Denna visas sedan i listrutan Urval när referensen infogas.  
I HTML-dokument tas dock ingen hänsyn till de referensfält som infogats på detta vis.  
Som mål för en korshänvisning i ett HTML-dokument måste Du infoga ett bokmärke.  
Infoga referens  
Infogar en korshänvisning till ett annat ställe i dokumentet.  
Det är bara då som Du kan infoga en hänvisning genom att välja ett fältnamn under Urval.  
I samlingsdokument kan Du även hänvisa från ett deldokument till ett annat.  
Här måste Du ta hänsyn till att referensens namn inte visas i urvalsfältet och att Du måste skriva in det "för hand".  
I HTML-dokument tas dock ingen hänsyn till de referensfält som infogats på detta vis.  
För korshänvisningar i HTML-dokument måste Du infoga en hyperlänk.  
Referenser är fältkommandon.  
Om du vill ta bort en referens raderar du fältkommandot.  
Sedan kan du infoga den igen som "oformaterad text" på samma ställe igen med kommandot Redigera - Klistra in innehåll.  
Då bibehålls själva texten medan referensen raderas.  
Om du har infogat ett bokmärke i dokumentet via Infoga - Bokmärke, så visas även posten "Bokmärken" under fliken Referenser.  
Bokmärken använder du för att markera vissa textavsnitt inom ett dokument.  
I ett textdokument kan du med hjälp av infogade bokmärken t.ex. snabbt hoppa från ett ställe i dokumentet till ett annat.  
I ett HTML-dokument förvandlas dessa bokmärken till ankare (A name) som t ex definierar hoppadressen för hyperlänkar.  
Namn  
Här skriver du in fältnamnet för nya fält som du definierar.  
Du tilldelar ett namn när du sätter en hoppadress.  
När du sedan infogar en referens till denna hoppadress, kan du identifiera hoppadressen med hjälp av namnet som visas i urvalsfältet för fälttypen "Sätt referens".  
När Du använder hänvisningar till ett samlingsdokuments olika deldokument, så måste Du skriva in namnet på en referens manuellt om den inte finns i samma deldokument.  
När Du sätter en referens till en markering i texten, så används den aktuella markeringen som fältinnehåll.  
Funktioner  
Här matar du in värden för fler funktionsparametrar.  
Typen av parametrar är beroende av den valda funktionen.  
Den kan vara kopplad till ett villkor beroende på fälttyp.  
Du kan definiera fält som utför ett visst makro när man klickar med musen, eller sådana som döljer textavsnitt om ett visst villkor uppfylls.  
För grafiska objekt, tabeller, ramar och andra objekt kan du definiera platshållare så att du kan infoga dem i dokumentet vid behov.  
Fälttyp  
Betydelse  
Villkorlig text  
Infogar en text om ett villkor uppfylls.  
Ange t.ex. "x eq 1" (utan citattecknen) under Villkor.  
Under Så skriver du en text som ska infogas i fallet x=1, och under Annars en text som infogas i övriga fall.  
X sätter du med fälttyperna "Sätt variabel" eller med ett inmatningsfält för en ny variabel (se Variabler).  
Inmatningsfält  
Infogar formulärfält för inmatning av text.  
Dessa kan Du förse med separata hänvisningar.  
När Du klickar på kommandoknappen Infoga, öppnas dialogrutan Inmatningsfält, där Du kan skriva in och redigera den önskade texten.  
Utför makro  
Infogar ett textfält som automatiskt utför ett tilldelat makro när du dubbelklickar.  
Du väljer det önskade makrot med kommandoknappen Makro....  
När du har valt makro skriver du in den tillhörande förklaringen i textfältet Hänvisning.  
Platshållare  
Infogar en platshållare i dokumentet.  
Platshållarens typ bestämmer Du under Format.  
Beteckningen skriver Du i textfältet Platshållare och eventuella förklaringar under Hänvisning.  
När Du klickar på platshållaren i dokumentet, kan Du infoga det objekt i vars ställe platshållaren står.  
Dold text  
Infogar en text som döljs om ett villkor är uppfyllt.  
Om du vill att sådana texter ska kunna döljas på bildskärmen, avmarkerar du rutan Dold text under Verktyg - Alternativ... - Textdokument - Formateringshjälp.  
Dolt stycke  
Döljer ett stycke om den förutsättning som du har registrerat under Villkor uppfylls.  
Det här fältkommandot kan du t.ex. använda så att tomma stycken döljs vid utskrift.  
Om du vill att sådana stycken ska döljas på bildskärmen, avmarkerar du menykommandot Visa - Dolda stycken eller kryssrutan Dolda stycken under Verktyg - Alternativ - Textdokument - Formateringshjälp.  
Villkoren för "Dold text" och "Dolt stycke "kan nu formuleras på samma sätt.  
StarWriter 4.0 gällde en omvänd logik för "Dold text".  
När du sparar och laddar äldre format, så omvänds därför logiken för "Dold text" automatiskt.  
Kombinera tecken (bara vid asiatiskt stöd)  
Här kan du kombinera 1 till 6 tecken som behandlas som ett standardtecken när kombinationen har gjorts.  
För funktionsfält används formatfältet bara för fältkommandon av typen platshållare.  
Här bestämmer du genom formatet för vilket objekt en platshållare gäller.  
Villkor  
Här anger du kriteriet för fält som är kopplade till ett villkor.  
Så, Annars  
Här kan Du ange fältinnehållen i relation till villkoret.  
Dessa tilldelas om villkoret är uppfyllt (Så) eller inte är uppfyllt (Annars).  
Dessa textfält är bara tillgängliga för funktionsfält av typen Villkorlig text.  
I resultatfälten Så och Annars kan du dels skriva in vanlig text, dels ange databasfält i form av "databasnamn.tabellnamn.fältnamn" (utan citattecken) så att fältinnehåll infogas om villkoret uppfylls. %PRODUCTNAME försöker vid sådana uttryck först identifiera texten som en databaskolumn.  
Om en sådan finns, så matas kolumnens innehåll ut, i annat fall bara texten.  
Om en villkorlig text innehåller ett uttryck med formen "databasnamn.databastabell.fältnamn" (utan citattecken), så tolkas den som databasuttryck och databasfältets tillhörande innehåll infogas.  
Ifall citattecknen sätts dit, så tolkas och infogas uttrycket som text.  
Citattecknen tas automatiskt bort innan fältinnehållet visas.  
Om det angivna tabell - eller fältnamnet inte finns i någon databas, så infogas ingenting om citattecknen inte sätts ut.  
Om det angivna databasnamnet inte motsvarar någon databas som är registrerad i %PRODUCTNAME, så tolkas och infogas uttrycket som text.  
Hänvisning  
Här anger du hänvisningen för respektive fälttyp.  
Urval  
Här väljer Du det makro som ska utföras ur en aktuell modul.  
Ifall den valda modulen bara innehåller ett makro, så finns också bara en post i urvalsfältet.  
Makronamn  
För fält som används för att köra ett makro visas här namnet på det makro som är markerat i urvalsfältet.  
Platshållare  
Här kan du definiera en platshållare när fälttypen Platshållare är vald.  
Infoga text  
När Du har valt fälttypen Dold text, kan Du skriva in den text som är kopplad till ett villkor här.  
Tecken  
Om du har valt fälttypen Kombinera tecken kan du ange tecknen som ska kombineras här.  
Värde  
Om du har valt fälttypen Kombinera tecken kan du ange ett värde här.  
Makro...  
Om du klickar på den här kommandoknappen öppnas dialogrutan Makro, där du kan välja ut ett makro som ska utföras när du klickar på fältkommandot.  
Den här kommandoknappen är bara aktiv om du har valt ett funktionsfält av typen "Utför makro".  
Dokumentinfo  
Dokumentinfofält innehåller data från dokumentegenskaperna.  
Till dessa hör dels allmänna uppgifter som %PRODUCTNAME automatiskt genererar och förvaltar för varje dokument, t.ex. data om när dokumentet har skapats och ändrats, dels manuellt inmatad information som du kan definiera individuellt för dokumentet.  
Innehållet i dokumentinfofälten är arkiverade i %PRODUCTNAME under Arkiv - Egenskaper.  
När dokumentinfofält importeras och exporteras i HTML-format, gäller speciella %PRODUCTNAME -format.  
Fälttyp  
Betydelse  
Ändring  
Infogar författarnamn, datum och / eller klockslag för den senaste gången som dokumentet sparades.  
Redigeringstid  
Infogar den tid som dokumentet redan har redigerats.  
Beskrivning  
Infogar dokumentbeskrivningen om denna har registrerats i dokumentegenskaperna.  
Dokumentnummer  
Infogar det aktuella dokumentnumret.  
Skapad  
Infogar författarnamn, datum och / eller klockslaget då dokumentets skapades.  
Info 0 - 3  
Infogar innehållet i dokumentegenskapernas infofält.  
Under Arkiv - Egenskaper... - Användare kan Du redigera infofältens innehåll.  
Senaste utskrift  
Infogar datum och / eller klockslag och / eller författarnamn för senaste utskriften.  
Nyckelord  
Infogar de nyckelord som har registrerats under Arkiv - Egenskaper... - Beskrivning.  
Tema  
Infogar det tema som har registrerats i dokumentegenskaperna.  
Rubrik  
Infogar den rubrik som har registrerats i dokumentegenskaperna.  
För dokumentinfofält kan Du välja mellan fältkommandona Författare, Klockslag och Datum när Du vill infoga fält av typen Ändring, Skapad och Senaste utskrift.  
Här kan Du ställa in datum - och tidformat för de aktuella fälttyperna.  
Fixera innehåll  
Om du har markerat den här rutan, så tilldelas fältet bara ett innehåll när det infogas i dokumentet och ändras sedan inte mer.  
Fält vars innehåll är fixerat tolkas alltid på nytt om ett nytt dokument skapas från en mall eller om ett textblock med ett fixerat fält infogas.  
Liksom med datumfälten används de data som gäller när dokumentet skapas från mallen eller när textblocket infogas.  
På så sätt säkerställs att globala mallar och textblock kan användas individuellt.  
Textblock med sådana fält kan Du t ex använda för signaturer.  
Variabler  
Med variabelfält styr du dokumentets innehåll dynamiskt.  
Du kan definiera variabler individuellt eller välja dem bland förinställda variabeltyper.  
Användardefinierade fält är bara tillgängliga i det aktuella dokumentet.  
Fälttyp  
Betydelse  
Sätt variabel  
Definition av en variabel och inmatning av variabelvärdet.  
Du kan ändra värdet på en definierad variabel med hjälp av inmatningsfältet, så att variabeln får olika värden på olika ställen i dokumentet.  
Visa variabel  
Infogar en variabels aktuella värde.  
Om Du har definierat en variabel med fälttypen "Sätt variabel" eller ändrat dess värde med fälttypen "Inmatningsfält", så kan Du infoga variabelns aktuella värde i dokumentet med ett fält av typen "Visa variabel ".  
Det aktuella variabelvärdet i dokumentet bestäms av föregående fält av typen "Sätt variabel" eller av det föregående inmatningsfältet.  
DDE-fält  
Infogar en DDE -länk som Du kan infoga i dokumentet och uppdatera så ofta Du vill via det fältnamn som Du har definierat.  
Infoga formel  
Infogar beräkningar eller fasta siffervärden.  
Du väljer önskat talformat under Format.  
Inmatningsfält  
Infogar ett nytt värde för en redan definierad variabel eller för ett användarfält.  
För ett inmatningsfält för en variabel gäller det nytilldelade värdet alltid från den position där Du infogar inmatningsfältet i dokumentet, och till dess att Du ändrar värdet genom att infoga ytterligare ett inmatningsfält.  
Vid ett inmatningsfält för ett användarfält ändrar Du användarfältets värde globalt, dvs det nya värdet gäller för varje användarfält i dokumentet.  
När du klickar på kommandoknappen Infoga, öppnas dialogrutan Inmatningsfält, där du kan skriva in det nya värdet tillsammans med en hänvisning.  
Nummersekvens  
Infogar en automatisk numrering för tabeller, grafiska objekt och textramar.  
Sätt sidvariabel  
Infogar en andra sidnumrering.  
Med "av" upphäver Du den.  
Visa sidvariabel  
Visar sidnumret, räknat från en referenspunkt.  
Du bestämmer referenspunkten med fälttypen "Sätt sidvariabel".  
Användarfält  
Individuell definition av en global variabel som t.ex. kan användas för att styra programhändelser.  
Du kan ändra ett användarfälts värde om du tilldelar användarfältet ett inmatningsfält.  
En ändring kan bara ske globalt och påverkar hela dokumentet.  
Om inte några användarfält är listade under Urval ännu, måste du först tilldela ett fältnamn och ett värde.  
Om du sedan klickar på ikonen Överta, så visas namnet på det användardefinierade fältet i urvalsfältet.  
För fält som Du definierar själv kan Du antingen välja det önskade formatet bland de förinställda formaten eller så klickar Du på posten "Ytterligare format..." för att bestämma ett eget format i dialogrutan Talformat.  
När det gäller nummersekvenser eller sidvariabler har du, utöver de vanliga numreringsformaten, även tillgång till numreringar med likadana små (a,... aa,... aaa) eller stora bokstäver (A,...  
AA,...  
AAA).  
I listrutan Format anger du om det registrerade värdet ska infogas i textformat eller i ett numeriskt format.  
I ett HTML-dokument har Du här för fälttypen "Sätt variabel" tillgång till fältkommandona HTML_ON och HTML_OFF.  
Dessa medför att den satta variabeln för HTML-källtexten konverteras till en inledande tagg (<Värde>) och en avslutande (< / Värde>), varvid posten under Värde infogas som text mellan vinkelparenteserna.  
Du kan även markera den önskade variabeln och trycka på blankstegstangenten.  
Formel  
Här anger Du formeln om Du har valt ett fält av typen "Infoga formel".  
Osynligt  
Om du markerar den här rutan, visas inte fältinnehållet i dokumentet.  
I stället för fältvärdet visas då bara en smal fältmarkering i dokumentet.  
Denna funktion är bara tillgänglig för de användardefinierade fälten "Sätt variabel" och Användarfält.  
Numrering kapitelvis  
I det här området anger du hur numreringen av kapitel ska börja om.  
Nivå  
Här väljer du den överskrifts - respektive kapitelnivå vid vilken numreringen ska börja om när nivån ändras.  
Skiljetecken  
Ange här det tecken som ska följa direkt efter numret på överskrifts - respektive kapitelnivå.  
Överta  
Med den här ikonen övertar du det användardefinierade fältkommandot till urvalslistan.  
Radera  
Med den här ikonen raderar du ett användardefinierat fältkommando från urvalslistan.  
Du kan bara radera fältkommandon om de inte finns i dokumentet.  
Om du har infogat ett fältkommando i dokumentet och vill ta bort den motsvarande posten från urvalslistan, så måste du först radera fältkommandot i dokumentet.  
Radera  
Databas  
Här kan du infoga databasfält från en databasfil.  
Bland fältkommandotyperna hittar du även standardbrevfält som du kan använda när du skapar standardbrev (kopplad utskrift).  
Vid kopplad utskrift infogar dessa fältkommandon fältinnehåll som är beroende av dataposterna.  
Fälttyp  
Betydelse  
Slumpvis datapost  
Om villkor et är uppfyllt, infogas innehållet i den datapost som du har definierat under Datapostnummer i ett efterföljande fält för kopplad utskrift.  
Hänsyn tas enbart till de dataposter som du har valt via en multimarkering i datakällvyn.  
Med hjälp av detta fältkommando kan Du infoga flera speciella dataposters innehåll på en dokumentsida.  
Då infogar Du ett fältkommando av typen Slumpvis datapost framför de fält för kopplad utskrift för vilka en viss datapost ska användas.  
Databasnamn  
Infogar namnet på den databasfil som Du kan välja i fältet till höger.  
Observera:  
Fältkommandot Databasnamn finns bara globalt.  
Ändrar Du något databasnamn, så ändras även alla andra i dokumentet.  
Datapostnummer  
Infogar numret på den datapost som är markerad.  
Välj den önskade formateringen under Format.  
Nästa datapost  
Om villkoret är uppfyllt, infogas innehållet i nästa datapost i ett efterföljande fält för kopplad utskrift.  
Hänsyn tas enbart till de dataposter som du har markerat via en multimarkering i datakällvyn.  
Med hjälp av detta fältkommando kan Du infoga innehållen för flera dataposter som följer efter varandra på en dokumentsida.  
Då infogar Du ett fältkommando av typen Nästa datapost mellan de fält för kopplad utskrift där ett byte av dataposten ska ske.  
Standardbrevfält  
Infogar namnet på ett databasfälts som platshållare.  
Fältinnehållet skrivs in automatiskt vid utskrift av standardbrev (kopplad utskrift).  
Databasurval  
Här kan Du välja en databastabell eller en sökning till vilken fältkommandot ska relatera.  
Du kan välja bland samtliga databaser som är registrerade i %PRODUCTNAME.  
På så vis kan Du integrera fältinnehållen från olika databaser, -tabeller eller -sökningar i ett dokument.  
Fält av typen "Slumpvis datapost" och "Nästa datapost "kan kopplas till ett villkor.  
Data i den angivna dataposten eller i nästa datapost infogas i dokumentet enbart om villkoret är uppfyllt.  
Villkoret är m a o alltid uppfyllt om Du inte ändrar villkorstexten.  
Datapostnummer  
Här anger du för fälttypen "Slumpvis datapost" datapostnumret på den datapost vars innehåll ska infogas om kriteriet under Villkor är uppfyllt.  
Datapostnumret relaterar alltid till den aktuella markeringen i datakällvyn.  
Det innebär t.ex. att om du i en databas med 10 dataposter bara har markerat de sista fem dataposterna, så väljer du med datapostnumret 1 den första markerade dataposten, d.v.s. den sjätte posten i den aktuella tabellen.  
Om du refererar till fälten i en annan databas (eller en annan tabell eller sökning inom samma databas), så bestäms datapostnumret relativt i förhållande till den aktuella markeringen.  
Om t.ex. en markering i den aktuella databastabellen inte omfattar den första dataposten, så innebär det att du med datapostnummer 1 inte anropar den första dataposten, utan den andra, i den andra databasen (eller i den andra tabellen eller sökningen).  
Format  
Här väljer Du det format i vilket fältinnehållet ska infogas.  
Dessa inställningar kan Du bara välja för datumfält.  
Från databas  
När Du väljer det här alternativet används formaten från databasen.  
Användardefinierat  
När Du väljer det här alternativet kan Du välja ett användardefinierat format från listan.  
Lista över användardefinierade format  
Här är alla användardefinierade format tillgängliga.  
Speciella taggar  
Här följer en förklaring av speciella taggar som används för fältkommandon.  
Om du skapar HTML-dokument med fältkommandon med hjälp av %PRODUCTNAME Writer, konverteras fältkommandona från %PRODUCTNAME till speciella taggar för HTML-källtexten.  
Dessa taggar är inte definierade i HTML-format, eftersom de avser specifika funktioner i %PRODUCTNAME, i det här fallet fältkommandon.  
När du importerar och exporterar HTML-dokument måste du därför tänka på att %PRODUCTNAME har egna internt definierade format för fältkommandon.  
Taggen för ett fältkommando i %PRODUCTNAME Writer är SDFIELD.  
Starttaggen innehåller alternativ för att ange fälttyp, format och det speciella fältet.  
Formatet för en fältkommandotagg, som känns igen av HTML-filtret, beror på fältkommandot.  
Dokumentfält av typen datum eller klockslag  
För dokumentfälten Datum och Klockslag anger Du DATETIME som värde för TYPE-alternativet.  
Alternativet SDNUM anger fältformatet, där det görs åtskillnad mellan datum - och klockslagsfält med hjälp av det där angivna formatet (t ex DD:MM:ÅÅ eller HH:MM:SS).  
Vid fasta datum - och klockslagsfält anger Du datum respektive klockslag med alternativet SDVAL.  
Det här alternativet avgör också om fältet är fast eller inte.  
I följande tabell kan Du med hjälp av exempel se vilka format för datum - respektive klockslagsfält som tolkas rätt av HTML-filtret:  
Fältkommando  
%PRODUCTNAME -tagg  
Datum fast  
<SDFIELD TYPE=DATETIME SDVAL=" 35843,4239988426 "SDNUM="1031;1031;DD.MM.ÅÅ ">17.02.98< / SDFIELD>  
Datum variabel  
<SDFIELD TYPE=DATETIME SDVAL=" 35843,4239988426 "SDNUM="1031;1031;DD.MM.ÅÅ ">17.02.98< / SDFIELD>  
Klockslag fast  
<SDFIELD TYPE=DATETIME SDVAL=" 35843,4240335648 "SDNUM="1031;1031;HH:MM:SS ">10:10:36< / SDFIELD>  
Klockslag variabelt  
<SDFIELD TYPE=DATETIME SDVAL=" 35843,4240335648 "SDNUM="1031;1031;HH:MM:SS ">10:10:36< / SDFIELD>  
Det gamla formatet stöds fortsättningsvis vid import.  
Det innebär m a o att Du inte längre kan skapa några fält som motsvarar äldre Office-versioner.  
Exempel för 4.0-formatet:  
<SDFIELD TYPE=DATE FORMAT=SSYS VALUE=" 19980217 ">17.02.98< / SDFIELD>  
<SDFIELD TYPE=TIME FORMAT=SYS VALUE=" 10083682 ">10:08:36< / SDFIELD>  
Dokumentinfofält  
För dokumentinfofälten anger du DOCINFO som värde för alternativet TYPE.  
Alternativet SUBTYPE anger den speciella fälttypen.  
Fältet av typen Skapa har SUBTYPE-alternativet CREATE, fälttypen Ändring har alternativet CHANGE.  
Formatet för dessa fält anges med alternativet SDNUM.  
Dessutom finns alternativet SDFIXED, som talar om att innehållet i dokumentinfofältet är fast.  
Om ett fast fält inte beskriver något datum eller klockslag, används texten mellan öppningstaggen <SDFIELD> och stopptaggen < / SDFIELD> som innehåll i fältet.  
Vid datum - och klockslagsfält anges fältets värde i ett SDVAL-alternativ.  
Exempel:  
Fältkommando  
%PRODUCTNAME -tagg  
Beskrivning (innehåll fast)  
<SDFIELD TYPE=DOCINFO SUBTYPE=COMMENT SDFIXED>beskrivning< / SDFIELD>  
Skapande datum  
<SDFIELD TYPE=DOCINFO SUBTYPE=CREATE FORMAT=DATE SDNUM=" 1031;1031;KK ÅÅ ">1 kvartalet 98< / SDFIELD>  
Skapande klockslag (innehåll fast)  
<SDFIELD TYPE=DOCINFO SUBTYPE=CREATE FORMAT=TIME SDVAL=" 0 "SDNUM="1031;1031;HH:MM:SS AM / PM" SDFIXED>03:58:35 PM< / SDFIELD>  
Ändring datum  
<SDFIELD TYPE=DOCINFO SUBTYPE=CHANGE FORMAT=DATE SDNUM=" 1031;1031;NN DD.MMM ÅÅ ">Må 23 feb 98< / SDFIELD>  
Inmatningsfält  
I den här dialogrutan definierar Du ett inmatningsfält.  
Det finns två typer av inmatningsfält, som kan infogas i dokumentet:  
Funktionsfält av typen inmatningsfält använder Du för textinmatning, medan Du använder variabelfält av typen inmatningsfält för att definiera nya variabelvärden.  
Om Du träffar på ett fältkommando av typen inmatningsfält i ett dokument, växlar pekaren utseende till en hand med utsträckt pekfinger.  
Om Du klickar öppnas den här dialogrutan, och Du kan redigera den text eller det värde som visas i det nedre textfältet.  
Redigera  
I det nedre textfältet anger Du den text eller det värde som ska visas.  
Nästa  
Genom att klicka på den här kommandoknappen går du till nästa inmatningsfält i dokumentet.  
Den här kommandoknappen visas bara om du har placerat markören framför ett inmatningsfält och tryckt på tangentkombination Skift+Ctrl+F9.  
Formulering av villkor  
Det finns kommandon som är kopplade till ett villkor, så att du kan styra utmatningen av dokumentinnehåll.  
I %PRODUCTNAME Writer formuleras i huvudsak villkor för fältkommandon, men det går även att göra visningen av definierade områden beroende av ett villkor.  
Men de här förklaringarna kan även tillämpas på områden.  
Villkor är nämligen logiska uttryck vars syntax, oberoende av sammanhanget, alltid är densamma i %PRODUCTNAME Writer.  
För fältkommandon kan du formulera villkor för följande fälttyper:  
Villkorlig text:  
Den infogade texten är kopplad till ett villkor.  
Om villkoret är sant infogas text A, i annat fall infogas text B.  
Dold text:  
Den infogade texten döljs om ett villkor är sant.  
Dolt stycke:  
Ett stycke i dokumentet döljs om ett villkor är sant.  
Slumpvis och Nästa datapost:  
Villkor i dessa databasfält styr åtkomsten till data som ska infogas i dokumentet ur en eller flera databaser.  
Du måste av princip alltid skriva in ett logiskt uttryck som villkor, eftersom ett villkor alltid är sant (uppfyllt) eller falskt (inte uppfyllt).  
Om ett logiskt uttryck är falskt så får det i %PRODUCTNAME värdet 0 (False), ifall uttrycket är sant så är värdet inte lika med 0 (True).  
Den enklaste sättet att ange en villkorstext är därför att direkt ange ett värde:  
True  
Villkoret är alltid uppfyllt.  
Du kan även ange ett valfritt värde inte lika med 0 som villkorstext.  
False  
Villkoret är inte uppfyllt.  
Du kan även ange värdet 0.  
Ett tomt villkorsfält tolkas som om villkoret inte är uppfyllt.  
Om textfältet Villkor är tomt, så ger det samma resultat som när du anger False eller 0.  
När du formulerar ett villkor kan du använda samma element som finns i formellisten när du formulerar en formel: operatorer, matematiska och statistiska funktioner, talformat, variabler och konstanter.  
De jämförande och logiska operatorerna är de grundläggande elementen som du behöver för att kunna formulera ett villkor.  
När du formulerar villkor kan du använda följande variabler:  
Användardefinierade variabler (fältkommando "Sätt variabel "eller Användarfält)  
Fördefinierade variabler i %PRODUCTNAME som tar upp statistiska värden ur dokumentegenskaperna  
Användardata  
Innehåll i databasfält  
Du kan dock inte använda de interna variablerna (sidnummer, kapitel osv) för ett villkor.  
Villkor och variabler  
X kan antingen vara namnet på ett egendefinierat fältkommando ("Sätt variabel "eller Användarfält) med ett definierat värde eller en %PRODUCTNAME -variabel vars värde är beroende av dokumentet.  
Exempel:  
x == 1 eller x EQ 1  
Villkoret är sant om variabeln x är lika med 1.  
Om Du exempelvis vill formulera ett villkor som tar hänsyn till det totala antalet sidor i dokumentet, så anger Du för x "Page":  
Page == 1 medför att villkoret blir sant om dokumentet bara innehåller en sida.  
x != 1 eller x NEQ 1  
Villkoret är sant om variabeln x inte är lika med 1.  
sinx == 0  
Villkoret är sant om variabeln x är en multipel av pi.  
Relationsoperatorer kan Du även använda för strängar.  
Dessa måste Du vanligtvis ange med dubbla citattecken:  
x == "ABC" eller x EQ "ABC "  
Kontrollerar om variabeln x innehåller strängen "ABC" (sant) eller inte (falskt).  
x == "" eller x EQ ""  
respektive  
!x eller NOT x  
Kontrollerar om variabeln x innehåller en tom sträng.  
Här övertar båda möjligheterna samma funktion.  
Du måste sätta två likhetstecken i villkoret för den jämförande operatorn "Lika med", t.ex. x == 1.  
Om du t.ex. har definierat en variabel med värdet 1 och sedan anger x = 1 som villkor, kan %PRODUCTNAME inte tolka ditt villkor korrekt och returnerar alltid värdet Falskt som resultat.  
Användardata  
När du formulerar ett villkor har du också åtkomst till de användardata som finns under Verktyg - Alternativ - %PRODUCTNAME - Användardata.  
Användardata består alltid av strängar, och du kan kontrollera innehållet med "==" (EQ) eller "!= "(NEQ) eller" !"(NOT).  
Variablernas namn i användarinformationen definieras så här:  
Variabel  
Betydelse  
user_firstname  
Förnamn  
user_lastname  
Efternamn  
user_initials  
Initialer  
user_company  
Företag  
user_street  
Gata  
user_country  
Land  
user_zipcode  
Postnummer  
user_city  
Ort  
user_title  
Titel  
user_position  
Befattning  
user_tel_work  
Telefon - arbetet  
user_tel_home  
Telefon - privat  
user_fax  
Faxnummer  
user_email  
E-postadress  
user_state  
Stat (inte i alla %PRODUCTNAME -versioner)  
Då anger Du som villkor: user_initials==" LM ".  
Villkor och databasfält  
När Du arbetar med databaser, kan Du formulera villkor som anropar innehållen i databasfält.  
Du kan dels använda villkor som kontrollerar om ett databasfält har något innehåll, dels sådana med vilka Du hämtar innehållet i ett databasfält.  
Även här tolkas logiska uttryck som har formulerats med hjälp av jämförande eller logiska operatorer.  
Några exempel:  
Exempel  
Betydelse  
databas.tabell.företag  
respektive  
databas.tabell.företag != "" eller databas.tabell.företag NEQ ""  
Returnerar Sant om datafältet FÖRETAG är fyllt. (I den första varianten behövs ingen operator.)  
!databas.tabell.företag eller  
NOT databas.tabell.företag  
respektive  
databas.tabell.företag == "" eller databas.tabell.företag EQ ""  
Returnerar Sant om datafältet FÖRETAG är tomt. (Utropstecken betyder logiskt NOT.)  
databas.tabell.företag != "Sun Microsystems" eller databas.tabell.företag NEQ "Sun Microsystems "  
Returnerar Sant om det aktuella värdet för datafältet FÖRETAG inte lyder "Sun Microsystems".  
databas.tabell.förnamn AND databas.tabell.namn  
Returnerar Sant om dataposten innehåller både för - och efternamn.  
Observera skillnaden mellan det logiska Inte "!" (NOT) och relationsoperatorn Inte lika med "!= "(NEQ).  
Som Du redan kan se i de ovanstående exemplen, så anges databasfält i formen "databasnamn.tabellnamn.fältnamn" (utan citattecken). %PRODUCTNAME upptäcker då automatiskt att det rör sig om ett databasfält.  
Då tolkas den som "normal" text av programmet.  
Exempel: dolt stycke i ett databasfält  
Anta att du har infogat ett fält för kopplad utskrift, FÖRETAG, i ett dokument.  
Men din adressboksdatakälla innehåller dataposter i vilka fältet FÖRETAG är tomt och därför skapas ett tomt stycke i ditt dokument.  
Detta stycke ska inte visas om datafältet är tomt.  
Välj fältkommandot Dolt stycke och ange som villkor: adressbok.adresser.företag EQ "" eller NOT adressbok.adresser.företag.  
Om databasfältet FÖRETAG är tomt, så är villkoret sant och stycket döljs och ignoreras vid utskrift.  
Om du har markerat kryssrutan Verktyg - Alternativ - Textdokument - Formateringshjälp - Dolda stycken, visas de dolda styckena på bildskärmen igen.  
Exempel på villkor i fältkommandon  
För alla fältkommandon som är kopplade till ett villkor finns samma möjligheter att formulera villkor.  
Detta illustreras med hjälp av fältet Villkorlig text nedan.  
Du kan dock utan vidare överföra syntaxen för ett villkor till fälten Dold text, Dolt stycke, Slumpvis eller Nästa datapost.  
Villkorlig text med en %PRODUCTNAME -variabel  
Öppna ett tomt textdokument och infoga ett fältkommando av typen Villkorlig text med följande parametrar:  
Villkor: page == 1  
Så:  
Det finns bara en sida.  
Annars:  
Det finns flera sidor  
Infoga sedan en manuell sidbrytning (menyn Infoga - Manuell brytning...) och tryck på F9 för att uppdatera fältinnehållet.  
Villkorlig text med en egendefinierad variabel  
Välj det numeriska formatet "Valuta" och infoga fältkommandot i dokumentet.  
Infoga nu ett fältkommando av typen Villkorlig text med följande parametrar:  
Villkor:  
Vinst < 10000  
Så:  
Uppsatt mål har inte nåtts.  
Annars:  
Uppsatt mål har nåtts.  
Öppna dialogrutan för redigering av fältkommandon genom att dubbelklicka på variabelfältet och ändra värdet från 5000 till 15000.  
Om Du bekräftar med OK, innebär det att uppsatta målet har nåtts.  
Villkorlig text med ett databasfält  
Öppna en datakälla och visa dataposterna.  
Infoga de två fälten FÖRNAMN och NAMN för kopplad utskrift direkt efter varandra i dokumentet.  
Markera en datapost i datakällvyn och klicka på ikonen Data i fält.  
Den markerade datapostens fältinnehåll infogas i dokumentet.  
Om förnamn saknas, ska blanksteget inte infogas.  
Placera markören mellan de båda fältkommandona och infoga ett extra fältkommando av typen Villkorlig text med följande parametrar:  
Villkor: adressbok.adresser.förnamn  
Så:  
Blanksteg  
Annars: (inget)  
Blanksteget infogas om ett förnamn har registrerats i adressboken.  
Då ser du att enbart efternamnet infogas.  
Villkor som refererar till databasfält kan Du överta till textfältet genom att dra och släppa dem.  
Förutom att Du i villkor kan kontrollera om ett datafält är fyllt, kan Du även avläsa innehållet:  
Infoga ett fältkommando av typen Villkorlig text med följande parametrar:  
Villkor: adressbok.adresser.förnamn == "Michael"  
Så:  
Bäste  
Annars:  
Hej  
Gör ett mellanslag efter fältkommandot och infoga sedan förnamnet som fält för kopplad utskrift.  
Det finns en beskrivning av hur du skapar standardbrev (kopplad utskrift) här.  
Förteckningar  
Här finns undermenyer med vars hjälp du kan utföra följande: infoga en ny post i en förteckning, skapa och utforma olika förteckningar och infoga en post i en litteraturförteckning.  
Post...  
Förteckningar...  
Litteraturförteckningspost...  
Infoga förteckningspost  
Med den här funktionen öppnar du en dialogruta där du kan definiera den markerade texten som post i en förteckning.  
Det kan t.ex. röra sig om en innehållsförteckning, ett sakregister eller en användardefinierad förteckning.  
Om du vill ändra en införd förteckningspost i efterhand, placerar du markören på eller omedelbart framför den plats där du har infogat posten och väljer sedan Redigera - Förteckningspost....  
Om Du markerar kryssrutan Använd på alla liknande texter (se nedan), införs i förteckningen alla likadana textställen i den löpande texten.  
Däremot inkluderas inte de förekomster som finns i ramar, sidhuvuden, sidfötter eller bildtexter.  
Om Du vill att alla förekomster av en viss text ska inkluderas i förteckningen, kan Du göra en upprepad ökning i texten (med kommandoknappen Sök alla i dialogrutan Sök och ersätt markerar Du alla förekomster på en gång).  
Sedan ger Du menykommandot Infoga - Förteckningar - Post...  
Dialogrutan Infoga förteckningspost finns kvar på bildskärmen tills Du stänger den.  
Medan dialogrutan är öppen, kan Du markera flera ord i texten (genom att t ex placera markören där) och sedan klicka på OK.  
Det markerade ordet införs i förteckningen.  
Markering  
I det här området väljer Du förteckning och infogar en önskad post.  
Förteckning  
Här väljer Du i vilken förteckning den markerade texten ska visas som förteckningspost.  
Post  
Här skriver Du den text som ska visas i förteckningen.  
Enligt standardinställning står texten som är markerad i dokumentet här.  
Du kan ändra texten i det här fältet och på så vis lägga in poster som inte finns som text i dokumentet i förteckningen.  
Om Du pekar med muspekaren alldeles intill en sådan post, visas som tipshjälp namnet på förteckningen samt själva texten i posten.  
Om detta ska fungera måste Du dock ha aktiverat tipshjälpen eller den aktiva hjälpen på Hjälp -menyn.  
Sorteringskod 1  
Om Du vill skapa ett register där sakorden är uppställda på flera nivåer anger Du här "övertermen" på den högsta nivån, eller också väljer Du den "överterm "som det aktuella sakordet ska underordnas.  
Du kan t ex ange "Redigera" som första nyckelord ("överterm") och "markera allt "som underpost.  
I det färdiga registret visas då följande post alfabetiskt inordnad under R: "Redigera, markera allt".  
Sorteringskod 2  
Om Du vill skapa ett register där sakorden är uppställda på flera nivåer, anger Du här "övertermen" på nivå två, eller också väljer Du den "överterm "som det aktuella sakordet ska underordnas.  
Huvudpost  
Genom att markera det här alternativet för ett sakregister, anger Du att den aktuella texten ska vara en huvudpost.  
Sidnumret för den markerade texten formateras i sakregistret med ett annat format än sidnumren för de andra förekomsterna av samma text.  
Nivå  
Om Du så vill införs automatiskt poster med styckeformateringen "Rubrik X" (X = 1-10) i innehållsförteckningen.  
Posternas nivå motsvarar därvid rubriknivån.  
För en fritt definierad post kan Du här bestämma på vilken nivå den ska föras in.  
Den här funktionen kan Du bara använda för innehållsförteckningar och användardefinierade förteckningar.  
Använd på alla liknande texter  
Om den här kryssrutan är markerad, specialmarkeras alla de textställen i löptexten som är lika med den för tillfället markerade texten som förteckningsposter.  
Inte heller inkluderas text som står i ramar eller bildtexter i ramar.  
Om Du vill använda den här funktionen markerar Du först ett textavsnitt i dokumentet och öppnar sedan dialogrutan Infoga förteckningspost.  
Om Du däremot skriver in en post manuellt, kan Du inte låta likadana textavsnitt i dokumentet automatiskt föras in i förteckningen på detta sätt.  
Exakt sökning  
Bara hela ord  
Infoga  
Klicka här om Du vill skapa en ny förteckningspost eller bekräfta en ändring av en post som Du just redigerar.  
Du kan omedelbart fortsätta att skapa eller redigera en ny post.  
Stäng  
Klicka här för att stänga dialogen när Du är klar.  
Ny användardefinierad förteckning  
Med den här kommandoknappen öppnar Du dialogrutan Skapa ny användardefinierad förteckning.  
Namn  
Här anger Du namnet på en ny användardefinierad förteckning.  
Du kan sedan välja den som ny typ på fliken Förteckning.  
Infoga förteckning  
Här infogar du en förteckning vid markörens position i dokumentet.  
Det finns olika typer av förteckningar att välja på, och du kan definiera så många andra typer som du vill.  
Om markören står i en förteckning när du väljer menykommandot Infoga - Förteckningar - Förteckningar..., kan du redigera den aktuella förteckningen här.  
I dialogrutan visas en förhandsvisning av den valda förteckningstypen.  
Om du har tilldelat delar av förteckningen egna mallar, eller ändrat standardmallarna, finns de här ändringarna med i förhandsvisningen.  
Dialogrutan innehåller flera flikar.  
Om du väljer en annan förteckningstyp i listrutan Typ under fliken Förteckning, ändras i allmänhet utseendet på flikarna Förteckning, Poster och Mallar beroende på vilken typ du väljer.  
Här definierar du antalet kolumner för förteckningens innehåll.  
Förteckningens rubrik omfattar alltid en kolumn från vänster till höger marginal, såvida du inte infogar hela förteckningen på en flerkolumnig sida.  
Mallar  
Här definierar du vilka styckeformatmallar som ska användas för förteckningsrubriker, skiljetecken och poster på de olika nivåerna.  
Dessutom kan du redigera styckeformatmallarna från den här dialogrutan.  
Tilldelning  
Om du vill formatera en förteckning kan du tilldela rubrik, skiljetecken och varje förteckningsnivå en annan styckeformatmall.  
Nivåer  
Markera här nivån för den förteckning, vars styckeformatmall Du vill ändra.  
Styckeformatmallar  
Markera här den styckeformatmall, som Du vill tilldela den markerade posten i den vänstra listan.  
Klicka sedan på Tilldela.  
<  
Den styckeformatmall som Du har markerat under Styckeformatmallar tilldelas den förteckningsnivå som Du har markerat under Nivåer.  
Standard  
Om Du har ändrat en tilldelning av en styckeformatmall återställs den för den markerade förteckningsnivån under Nivåer till standardtilldelningen (dvs den tilldelning som gäller när %PRODUCTNAME är nyinstallerat).  
Redigera  
Öppnar dialogrutan Styckeformatmall, där Du kan redigera den markerade styckeformatmallen.  
Förteckning  
När du skapar en ny förteckning, bestämmer du först typ av förteckning här.  
Om du vill kan du skapa flera användardefinierade förteckningar (t.ex. genom att ange en post med kommandot Infoga - Förteckningar - Post).  
Den här fliken ändrar utseende och funktion beroende på vilken typ som valts.  
Innehållsförteckning  
Sakregister  
Illustrationsförteckning  
Tabellförteckning  
Användardefinierad  
Objektförteckning  
Litteraturförteckning  
Förteckning  
Funktionen för fliken Förteckning, när Du har valt "Innehållsförteckning" som Typ.  
Typ och rubrik  
Välj typ och rubrik för förteckningen här.  
Typ  
I den här listrutan väljer du typ av förteckning.  
Beroende på vad du har valt ändras funktionerna under flikarna Förteckning, Poster och Mallar.  
Då kan du inte välja typ.  
Rubrik  
Här kan du ge den aktuella förteckningstypen en valfri rubrik.  
Rubriken visas som förteckningens överskrift i dokumentet.  
Skyddad mot manuella ändringar  
Om du markerar den här rutan, skyddar du innehållet i förteckningen som skapats i dokumentet mot ändringar.  
Manuella ändringar som du gör i en skapad förteckning går förlorade nästa gång som förteckningen uppdateras.  
Du kan bläddra med markören genom ett skyddat område om du markerar rutan Markör i skyddade områden - Tillåt under Verktyg - Alternativ - Textdokument - Formateringshjälp.  
Skapa förteckning för  
Här väljer du om förteckningen ska skapas för hela dokumentet eller bara för det aktuella kapitlet.  
Utvärdera till nivå  
För en innehållsförteckning väljer Du här på vilken överskriftsnivå överskrifterna och de poster Du klassat i förteckningen ska visas.  
Skapa från  
I det här området definierar Du vilken information som ska sammanfattas till en förteckning.  
Om Du markerar flera kryssrutor, övertas alla markerade poster i förteckningen.  
Disposition  
Om Du markerar den här rutan, övertas de stycken i innehållsförteckningen som är aktiva för dispositionen av dokumentet.  
Det gäller stycken med mallarna "Överskrift 1" till "10 "och mallarna som används för kapitelnumrering.  
...  
Här kan du definiera vilka styckeformatmallar som ska gälla för de olika nivåerna i dispositionen.  
Ytterligare mallar  
Om du klickar på den här rutan, tas alla texter som försetts med vissa styckeformatmallar med i förteckningen.  
Mallarna och deras nivå i förteckningen definierar du i dialogrutan Tilldela mall, som du öppnar genom att klicka på kommandoknappen... efter rutan.  
...  
Öppnar dialogrutan Tilldela mall.  
Förteckningsmarkeringar  
Om du markerar den här rutan, beaktas alla poster som du har infogat som poster för förteckningen med menykommandot Infoga - Förteckningar - Post när du skapade förteckningen.  
Förteckning  
Funktionen för fliken Förteckning, när Du har valt "Sakregister" som Typ.  
Tillägg  
Med de här kryssrutorna påverkar Du sakregistrets uppbyggnad.  
Kombinera likadana poster  
Om sakregistret innehåller flera likalydande begrepp, sammanfattar %PRODUCTNAME begreppen enligt följande: "Visning 10, visning 43" blir till "visning 10, 43 ", varvid siffrorna avser sidnumren.  
Kombinera med f eller ff  
Om sakregistret innehåller flera identiska poster på sidor som följer på varandra, sammanfattar %PRODUCTNAME posterna enligt följande: "Visning 10, visning 11, visning 12" blir till "visning 10ff ".  
Enkelt "f" betyder en följande sida, "ff "betyder flera följande sidor.  
Kombinera med -  
Om sakregistret innehåller flera identiska poster på sidor som följer på varandra, sammanfattar %PRODUCTNAME posterna enligt följande: "Visning 10, visning 11, visning 12" blir till "visning 10-12 ".  
Observera stor och liten bokstav  
Markera den här kryssrutan, om poster med stor respektive liten begynnelsebokstav ska föras in separat i sakregistret.  
Den här kryssrutan är bara relevant, om likadana poster ska kombineras:  
Om Du markerar kryssrutan Kombinera likadana poster, sammanfattar programmet likalydande poster oavsett stor eller liten bokstav.  
Då bestämmer den första posten som påträffas i dokumentet, om posten ska skrivas med liten eller stor bokstav.  
Skriv automatiskt poster med stor bokstav  
Om Du markerar den här rutan, kommer alla poster i förteckningen som börjar med en bokstav att visas med stor bokstav.  
Nyckel som egen post  
Markera den här kryssrutan, om Du vill infoga ett nyckelbegrepp som egen post i förteckningen.  
De tilldelade begreppen placeras under nyckelordet med indrag.  
Du definierar nyckelbegrepp i dialogrutan Infoga förteckningspost.  
Konkordansfil  
Om du markerar den här rutan, tas hänsyn till konkordansfilen (överensstämmelsefilen) när sakregistret skapas.  
Fil  
Den här kommandoknappen visar en undermeny med kommandona Öppna, Ny... och Redigera...  
Öppna  
Visar dialogrutan Öppna, där du kan välja konkordansfil.  
Om konkordansfilen inte har tillägget *.sdi utan exempelvis *.txt, skriver du in *.txt i fältet filnamn.  
Då visas filerna med detta filnamnstillägg.  
Ny...  
Dialogrutan Spara som visas, där Du kan välja sökväg och filnamn för den konkordansfil som ska skapas.  
Välj helst filnamnstillägget *.sdi, eftersom denna filtyp visas först när Du öppnar dialogrutan vid senare tillfälle.  
Filen sparas som ren textfil utan formateringar.  
Om Du avslutade dialogrutan med Spara, visas dialogrutan Redigera konkordansfil.  
Redigera...  
Här öppnar Du dialogrutan Redigera konkordansfil.  
Sortera  
Definiera här på vilket sätt förteckningsposterna ska sorteras.  
Språk  
Välj språket för sorteringen här.  
Nyckeltyp  
Välj nyckeltypen för sorteringen här.  
Förteckning  
Funktionen för fliken Förteckning, när Du har valt "Illustrationsförteckning" som Typ.  
Skapa från  
I det här området definierar Du vilken information som ska sammanfattas till en förteckning.  
Bildtexter  
Om Du har markerat det här alternativet, skapas posterna i illustrationsförteckningen från bildtexterna.  
Du kan tilldela ett markerat objekt en bildtext med kommandot Infoga - Bildtext....  
Kategori  
Välj här den kategori, varifrån alla funna objekt ska läggs till i den aktuella förteckningen.  
När Du ger objekten bildtexter kan Du definiera egna nummersekvenser och välja en av dem som kategori.  
Visning  
Välj här vad som ska visas som post.  
I följande tabell visas de olika alternativen.  
Bildtexten lyder i det här exemplet: "Illustration 24:  
Solen". "Illustration 24 "har genererats automatiskt, och":  
Solen "har Du lagt till.  
Val i listrutan Visning  
Post i förteckningen  
Referenstext  
Illustration 24:  
Solen  
Kategori och nummer  
Illustration 24  
Bildtext  
Solen  
När Du väljer "Bildtext" tas skiljetecknet och blanksteget i början av Din egen text automatiskt bort.  
Objektnamn  
Med det här alternativet skapar du förteckningsposter av objektnamnen.  
Du kan t.ex. visa objektnamnen i Navigator och ändra där i snabbmenyn.  
Förteckning  
Funktionen för fliken Förteckning, när Du har valt "Tabellförteckning" som Typ.  
Förteckning  
Funktionen för fliken Förteckning, när Du har valt "Användardefinierad" som Typ.  
Den användardefinierade förteckningen med den förinställda typen "Användardefinierad" är bara en av alla de förteckningar som du kan definiera själv.  
Om du definierar en förteckningspost, kan du ange i vilken förteckning du vill ha den.  
I samband med detta kan du också definiera en egen förteckning och ge den en typ med eget namn.  
De förteckningar vars typ Du själv har definierat finns med och kan väljas som posten "Användardefinierad" i listrutan Typ på fliken Förteckning.  
Skapa från  
I det här området definierar du vilken information som ska sammanfattas till en förteckning.  
Mallar  
Tabeller  
Markera här om alla tabeller ska tas med i förteckningen.  
Grafik  
Markera här om alla grafiska objekt ska tas med i förteckningen.  
Textramar  
Markera här om alla textramar ska tas med i förteckningen.  
OLE-objekt  
Markera den här rutan om alla OLE-objekt ska tas med i förteckningen.  
Nivå från ursprungskapitel  
Om Du markerar den här rutan, dras posterna i tabellerna, grafikobjekten, textramarna och OLE-objekten i förteckningen in så långt som motsvarar den hierarkiska indragningen för kapitlets överskrift.  
Om rutan inte är markerad, visas alla funna poster på den första nivån.  
Förteckning  
Funktionen för fliken Förteckning, när Du har valt "Objektförteckning" som Typ.  
Skapa utifrån följande objekt  
Markera alla objekttyper som ska tas med i objektförteckningen i listrutan.  
Förteckning  
Funktionen för fliken Förteckning, när Du har valt "Litteraturförteckning" som Typ.  
Formatering av poster  
Här fastställer Du hur litteraturförteckningsposterna ska se ut i löptexten respektive förteckningen.  
Numrera poster  
Om Du markerar den här rutan, numreras litteraturförteckningsposterna löpande.  
Parenteser  
Här kan Du välja stil för litteraturhänvisningarnas parenteser.  
Tilldela mall  
Här tilldelar Du de styckeformatmallar som finns i dokumentet en nivå i förteckningen.  
Mallar  
I den stora listrutan visas alla styckeformatmallar som finns i dokumentet. (Det är inte nödvändigt att tilldela mallarna ett stycke - det räcker om Du dubbelklickar på flera mallar efter varandra i Stylist för att de ska föras in i den stora listrutan.)  
Först står alla mallar på vänster sida i kolumnen "Inte tilldelat".  
Markera en mall.  
Med kommandoknappen >> kan Du flytta den här mallen till någon av kolumnerna 1 till 10.  
Därigenom läggs all text som är formaterad med den markerade styckeformatmallen till en förteckning på den nivå i hierarkin som motsvarar kolumnnumret.  
<<  
Här placerar Du den markerade mallen en kolumn längre åt vänster.  
>>  
Här placerar Du den markerade mallen en kolumn längre åt höger.  
Poster (förteckningar)  
Här gör du inställningar av formatet för förteckningsposter.  
Beroende på vad du väljer under fliken Förteckning ändras funktionen under fliken Poster.  
Välj en förteckningstyp för mer information.  
Innehållsförteckning  
Sakregister  
Illustrationsförteckning  
Tabellförteckning  
Användardefinierad  
Objektförteckning  
Litteraturförteckning  
Poster (innehållsförteckning)  
Här gör du inställningar av posternas format i en innehållsförteckning.  
Nivå  
I området Struktur definierar du sedan hur en post i förteckningen ska vara uppbyggd för den här nivån.  
För innehållsförteckningar finns det 10 tillgängliga poster.  
Med posten 1-10 väljer Du en gemensam struktur och formatering för alla 10 nivåer.  
Struktur  
På strukturraden definierar du med hjälp av olika fält utseendet på de olika posterna i förteckningen.  
Tomma fält och fält med beteckningar visas omväxlande.  
Du kan klicka på ett tomt fält och skriva in valfri text.  
Egenskaperna för ett markerat fält ställer du in med de andra styrfunktionerna i området Struktur.  
Om raden blir för lång kan Du flytta visningen av strukturraden åt vänster eller höger med två knappar.  
Du raderar en förkortning genom att markera den och trycka på tangenten Delete.  
Du skriver över en förkortning med en annan förkortning genom att markera den och sedan klicka på kommandoknappen för den andra förkortningen.  
På strukturraden infogar du fler förkortningar genom att sätta markören i ett tomt fält och klicka på kommandoknappen för en förkortning.  
Följande förkortningar är tillgängliga:  
Kapitelnr  
Infogar hänvisningens kapitelnummer (E#).  
Posttext  
Infogar hänvisningens text (ET eller E).  
Tabulator  
Infogar en tabb (T).  
Sidnr  
Infogar hänvisningens sidnummer (#).  
Hyperlänk  
Infogar omväxlande förkortningen för en hyperlänks början (LS) respektive slut (LE).  
När du klickar på hyperlänken hoppar markören och visningen till målet i dokumentet.  
Du kan välja stycken som mål vars styckeformatmall är angiven under Verktyg - Kapitelnumrerng  
Alla nivåer  
Om Du klickar på den här kommandoknappen, övertas den aktuella nivåns inställningar på alla nivåer.  
Teckenformatmall  
Här kan Du välja en teckenformatmall för det fält som har markerats på strukturraden.  
Redigera  
Med den här kommandoknappen öppnar du en dialogruta, där du kan redigera den markerade teckenformatmallen.  
Det skapas alltså inte någon kopia eller ny formatmall.  
Utfyllnadstecken  
Här markerar Du i listan, eller skriver in, det utfyllnadstecken som ska placeras framför tabbpositionen.  
Tabulatorposition  
Definiera här tabbens position i förhållande till vänstermarginalen.  
Vid högermarginalen  
Om du klickar i den här rutan, högerjusteras tabben vid höger textmarginal.  
Formatering  
Här definierar du fler formateringar för posterna.  
Tabbarnas position relativ till indraget från styckeformatmallen  
Om du markerar den här rutan, gäller de angivna tabbpositionerna relativt i förhållande till "indraget från vänster" i den valda styckeformatmallen.  
Annars gäller de relativt i förhållande till vänster textmarginal.  
Poster (sakregister)  
Här gör du inställningar av posternas format i ett sakregister.  
Den första nivån med namnet T skiljer sig från de andra nivåerna: den avser endast skiljetecknen.  
Om Du har bockmarkerat Alfabetiskt skiljetecken i området Formatering, visas en egen rad med begynnelsebokstaven för de följande posterna.  
På nivå T definierar Du hur denna rad formateras varje gång.  
Kapitelinfo  
Infogar kapitelinformationen (CI).  
Om Du markerar en post av denna typ på strukturraden, och enbart då, visas listrutan Kapitelpost längre ned i området Struktur.  
Kapitelpost  
Markera här det som Du vill ska visas som kapitelinformation:  
Nummersekvens och beskrivning, Bara nummersekvens, Bara beskrivning.  
Teckenformatmall för huvudposter  
Här anger Du teckenformatmallen för huvudposterna i sakregistret.  
Att en hänvisning ska vara en huvudpost anger Du i dialogrutan Infoga förteckningspost.  
Alfabetiskt skiljetecken  
Markera den här rutan, om Du vill skapa en egen rad med begynnelsebokstaven för de följande posterna.  
Nyckel, kommaseparerad  
Om Du markerar den här rutan, visas inte posterna i förteckningen på var sin rad utan efter varandra, separerade med kommatecken.  
Poster (illustrationsförteckning)  
Här gör du inställningar av posternas format i en illustrationsförteckning.  
För illustrationsförteckningar finns bara Nivå 1.  
Poster (tabellförteckning)  
Här gör du inställningar av posternas format i en tabellförteckning.  
För tabellförteckningar finns bara Nivå 1.  
Poster (användardefinierad förteckning)  
Här gör du inställningar av posternas format i en användardefinierad förteckning.  
För användardefinierade förteckningar finns bara Nivå 1.  
Poster (objektförteckning)  
Här gör du inställningar av posternas format i en objektförteckning.  
För objektförteckningar finns bara Nivå 1.  
Poster (litteraturförteckning)  
Här gör du inställningar av posternas format i en litteraturförteckning.  
Som nivåer visas här litteraturhänvisningarnas olika källor.  
Beroende på källa anges vanligtvis andra rader i litteraturförteckningen:  
För tidskriftsartiklar måste t ex månaden anges, vilket inte är brukligt för böcker.  
Postdata  
I den här listrutan visas de data som Du kan ange i dialogrutan Definiera litteraturpost.  
Sätt markören i ett ledigt fält på strukturraden, välj ut en rad från listrutan och klicka på kommandoknappen Infoga.  
Infoga  
Sätt markören i ett ledigt fält på strukturraden, välj ut en rad från listrutan och klicka på kommandoknappen Infoga.  
Ta bort  
Sätt markören på en beteckning på strukturraden och klicka på kommandoknappen Ta bort, om Du vill ta bort beteckningen.  
Sortering efter...  
Ange här vad posterna i litteraturförteckningen ska sorteras efter.  
Dokumentposition  
Posterna i litteraturförteckningen sorteras efter hänvisningarnas position i dokumentet.  
Detta är särskilt meningsfullt om hänvisningarna numreras automatiskt.  
Innehåll  
Posterna i litteraturförteckningen sorteras efter innehåll, t ex efter författare och utgivningsår.  
Sorteringsnyckel  
Om Du har markerat "Sortering efter innehåll", kan Du ange sorteringsnyckeln här.  
1, 2 eller 3  
Välj sorteringsnyckeln från tillgängliga postdata här.  
AZ  
Klicka på den här symbolen, om Du vill göra en alfanumerisk stigande sortering.  
ZA  
Klicka på den här symbolen, om Du vill göra en alfanumerisk fallande sortering.  
Definiera litteraturpost  
Här definierar Du en posts egenskaper för en litteraturförteckning.  
Postdata  
Skriv in en kort beteckning här och välj en passande typ.  
Nu kan Du skriva in data som hör till den här posten i de andra fälten.  
Vilka av dessa data som ska visas i litteraturförteckningen, bestämmer Du på strukturraden på fliken Poster i dialogrutan Infoga förteckning.  
Kort beteckning  
Här anger Du den korta beteckningen.  
Välj data för din litteraturförteckning här.  
Typ  
Välj här typ av litteraturförteckningspost i listan.  
Fälten i litteraturdatabasen har följande namn:  
"Identifier"; "BibliographyType"; "Author"; "Title"; "Year"; "ISBN"; "Booktitle"; "Chapter"; "Edition"; "Editor"; "Howpublished"; "Institution"; "Journal"; "Month"; "Note"; "Annote"; "Number"; "Organizations"; "Pages"; "Publisher"; "Address"; "School"; "Series" ;"ReportType"; "Volume"; "URL"; "Custom1"; "Custom2"; "Custom3"; "Custom4"; "Custom5";  
Redigera konkordansfil  
I den här dialogrutan skriver Du in sakregisterposter radvis.  
Du öppnar dialogrutan med menykommandotInfoga - Förteckningar - Förteckningar... - fliken Förteckning - markera "Sakregister" - markera Konkordansfil - kommandoknappen Fil - menykommandot Nytt.. eller Redigera...  
"Sökbegrepp" är den text som påträffas i dokumentet.  
"Alternativpost" är den text som visas i förteckningen som post.  
Nycklarna 1 och 2 är överordnade poster, under vilka Du kan inordna posten om Du vill.  
"Exakt" betyder att versaler och gemener matchas.  
"Hela ord" betyder att sökbegreppet inte får vara del av ett ord utan är ett ord i sig.  
Bockmarkera alternativen "Exakt" och / eller "Hela ord", om Du vill sätta dem på "Ja ".  
Du kan även skapa en konkordansfil själv och spara den som "textfil" utan formatering, om Du inte vill använda dialogrutan Redigera konkordansfil.  
Följande format gäller:  
Varje post står på en egen rad i konkordansfilen.  
Rader som börjar med # gäller som kommentarer.  
Formatet för en post i konkordansfilen definieras enligt följande:  
Sökbegrepp; Alternativpost;1 nyckel;2 nyckel;Exakt ;Hela ord  
Posterna för "Exakt" och "Hela ord "tolkas som "Nej" eller FALSE, om de är 0 (siffran noll) eller tomma.  
Allt annat innehåll tolkas som "Ja" eller TRUE.  
Om Du t ex alltid vill ha med ordet Göteborg i sakregistret under posten "Städer", skriver Du in följande rad i konkordansfilen:  
Göteborg; Göteborg;Städer;;0 ;0  
Den här raden hittar Göteborg även med gemener eller som del av ett ord.  
Om Du även vill ta med stadsdelen Örgryte under det hierarkiska stickordet Städer som posten "Göteborg", infogar Du följande rad:  
Örgryte; Göteborg;Städer;  
Om Du vill visa Göteborg under den hierarkiska posten Sverige / Städer, blir raden så här:  
Göteborg; Göteborg;Sverige ;Städer  
Infoga litteraturförteckningspost  
Här infogar du en post för litteraturförteckningen.  
Post  
I det här området definierar du posten.  
Från litteraturdatabas  
Markera det här alternativet, om Du vill välja posten från databasen "Bibliografi".  
Från dokumentinnehåll  
Välj det här alternativet om du vill markera posten bland de poster som redan finns i det aktuella dokumentet.  
En post i dokumentinnehållet kan vara likadan som en post i litteraturdatabasen.  
Posten i dokumentet har högre prioritet.  
När ett dokument med litteraturförteckningsposter sparas, sparas all information som hör till posterna automatiskt i ett dolt fältkommando.  
Det sker oberoende av om litteraturförteckningen skapades i dokumentet eller ej.  
Kort beteckning  
Välj här den korta beteckningen från litteraturdatabasen eller från posterna i det aktuella dokumentet.  
Författare, titel  
Här visas författare och titel för den korta beteckning som Du har valt, förutsatt att de redan är kända i litteraturdatabasen eller i det aktuella dokumentet.  
Infoga  
Klicka här om Du vill infoga hänvisningen i texten.  
Om Du har definierat en ny datapost med kommandoknappen Ny, måste Du absolut infoga denna även som post, annars går dataposten förlorad när Du stänger dokumentet.  
Stäng  
Stänger dialogrutan.  
Ny  
Öppnar dialogrutan Definiera litteraturpost med en tom inmatningsmask.  
Du kan definiera en ny datapost, som sparas i dokumentet, om Du också infogar en post för denna datapost.  
Om Du vill skapa en ny datapost i litteraturdatabasen, använder Du menykommandot Redigera - Litteraturdatabas.  
Redigera  
Öppnar dialogrutan Definiera litteraturpost, där Du kan redigera den aktuella dataposten.  
Information om att arbeta med litteraturförteckningsposter.  
Ram  
Med den här funktionen skapar eller redigerar du en ram, även med flera kolumner.  
Välj menykommandot Infoga - Ram så öppnas en dialog där du definierar en ram som infogas i det aktuella dokumentet.  
Kommandot Ram... visas bara i menyn Format om du har markerat en ram.  
Du kan även ändra en markerad ram med speciella kortkommandon.  
Om en ram med fast höjd innehåller mer text än vad som kan visas, kan Du rulla texten med hjälp av piltangenterna.  
Små röda pilar i textens början och slut anger att det finns mer text där.  
I förhandsvisningen i dialogrutan Format - Ram markeras referensområdet med en röd kvadrat och själva ramen med en grön.  
I förhandsvisningen visas också vilken effekt justeringen mot baslinje, rad och tecken har på ramar som har infogats "som tecken". "Baslinjen" är den linje på vilken alla radens tecken står; med "tecken "menas den höjd som omsluter alla radens tecken inklusive nedstaplar; och med "rad" menas den totala radhöjden inklusive alla objekt som är infogade som tecken.  
För ramar som är förankrade "till tecken" finns ytterligare ett referensområde, nämligen "tecken ".  
Detta motsvarar den blinkande textmarkörens streck när det står framför det tecken som har valts som ankare.  
Om Du väljer detta i lodrät riktning, kan Du förutom Överst, Nederst och Mitten även ställa in "Nedifrån" med ett fast avstånd.  
Exempelvis placeras en ram med "Vänster / Textområde i stycke samt Nedifrån 0 cm / Tecken" alltid vid vänster textkant på den rad som följer efter ankartecknet.  
Ikon på utrullningslisten Infoga på verktygslisten:  
Med ikonen Infoga ram manuellt ritar du snabbt upp en ram i dokumentet.  
Ändra ramar, grafiska objekt och objekt per tangentbord  
Här följer en kort beskrivning av hur Du på ett enkelt sätt kan ändra ramar, grafiska objekt och objekt med tangentbordet.  
Om en ram, ett grafisk objekt eller ett OLE-objekt är markerat eller om textmarkören blinkar i en ram, så kan Du ändra det markerade objektet med hjälp av piltangenterna.  
Om Du vill flytta objektet, så använder Du motsvarande piltangent tillsammans med Alternativ Alt -tangenten.  
Om Du vill ändra objektets storlek, så kan Du flytta den högra / nedre kanten med kortkommandot Kommando+Alternativ Ctrl+Alt och motsvarande piltangent.  
Om Du vill flytta den vänstra / övre kanten, håller Du dessutom skifttangenten nedtryckt.  
En sådan flyttning eller storleksändring gör Du utifrån de rastersteg som Du har angett under Verktyg - Alternativ... - Textdokument - Raster.  
När Du förflyttar ramar som är bundna till stycken begränsas Du därför till den högra / vänstra marginalen.  
För ramar som är bundna till tecken begränsas förflyttningen till överst / centrerad och underst.  
Infoga tabell  
Med den här funktionen kan du infoga en tabell i dokumentet.  
Om markören redan står i en tabell när du väljer kommandot, öppnas dialogrutan Tabellformat.  
Du kan även infoga en tabell från ett annat dokument med hjälp av urklippet.  
Då bevaras t.o.m. komplicerade formateringar som sammanslagna celler.  
Tomma rader av sammanfogade celler ger skapar vare sig blanksteg eller radbrytningar.  
Naturligtvis kan du också ge den nya tabellen intressanta formateringar och rama in kolumner och rader med enkla linjer.  
Om du vill formatera ett textavsnitt i dokumentet som texttabell, markerar du texten och klickar sedan på ikonen Infoga tabell på verktygslisten.  
Du kan också markera textavsnittet och sedan välja kommandot Verktyg - Text <-> Tabell, om du vill bestämma några av tabellens egenskaper i förväg i en dialogruta.  
När du infogar värden i en texttabell i %PRODUCTNAME Writer, formateras de automatiskt (t.ex. automatiskt igenkänning av datumvärden, tal, klockslag).  
Den här automatiska formateringen kan du stänga av i området Inmatning i tabeller i dialogrutan som du öppnar med Verktyg - Alternativ - Textdokument - Tabell.  
Namn  
I det här textfältet anger du namnet på den nya tabellen.  
Du kan också godta programmets standardförslag, då döps tabellen till TabellX (X är ett löpnummer).  
Tabellstorlek  
Här finns två rotationsfält, där du anger kolumn - och radantal för den nya tabellen.  
Kolumner  
Här väljer du antalet kolumner i tabellen.  
Rader  
Här väljer du antalet rader i tabellen.  
Alternativ  
I det här området definierar du egenskaper för tabellen som ska infogas.  
Jämför även menykommandona Format - Tabell - Textflöde och Verktyg - Alternativ - Textdokument - Tabell.  
Överskrift  
Om tabellens överskrift ska följa med till den nya sidan efter en sidbrytning, väljer du det här alternativet.  
Upprepa på varje sida  
Det här alternativet är bara tillgängligt bara om du har aktiverat alternativet Överskrift.  
Om du markerar den här rutan, upprepas överskriften i förekommande fall på varje sida.  
Dela inte tabell  
Om du väljer det här alternativet förhindrar du en eventuell delning av tabellen.  
Inramning  
Om du vill att tabellcellerna ska ramas in klickar du på den här rutan.  
Autoformat...  
Med den här kommandoknappen öppnar du dialogrutan Autoformat, där du kan välja layout för den nya tabellen.  
När du har stängt dialogrutan med OK, är du tillbaka i dialogrutan Infoga tabell, och den nya tabellen infogas med den valda layouten.  
Om du däremot klickar på Avbryt i dialogrutan AutoFormat, används ingen layout.  
Ikon på utrullningslisten Infoga på verktygslisten  
Om du väljer menykommandot Infoga - Tabell eller klickar kort på ikonen Tabell, öppnas dialogrutan Infoga tabell, där du definierar en tabell innan du infogar den i dokumentet med OK.  
När du släpper upp musknappen, infogas tabellen i dokumentet.  
Om det redan finns en tabell i dokumentet och markören står i den, öppnas dialogrutan Tabellformat när du klickar på ikonen.  
Det finns en begränsning för den maximala storleken på en tabellcell för närvarande: det får inte stå mer text i en cell än vad som får plats på en sida.  
Det är inte möjligt att göra en sidbrytning i en tabellcell.  
När du bläddrar genom ett textdokument med en tabellcell som är större än en sida hör du en varningssignal.  
Byt databas  
Här byter du ut databasen som du använder i det aktuella dokumentet mot en annan.  
Detta fungerar bara om databasfälten som du har infogat i dokumentet har samma fältnamn i båda databaserna.  
Om Du t ex har definierat en kopplad utskrift med adressfält från en databas men nu vill skicka utskriften även till mottagarna i databas B, behöver Du inte ersätta alla infogade fält utan bara byta databaser.  
De datafält i databas A som Du har infört i dokumentet ersätts av datafälten med samma namn i databas B.  
Observera informationen längre fram i detta avsnitt.  
Byt databas  
Du kan bara göra en sådan ändring per arbetspass.  
Använda databaser  
I den här listrutan visas vilka databaser som används i dokumentet.  
Från varje databas i listan har minst ett datafält infogats i dokumentet.  
Tillgängliga databaser  
I den här listrutan visas alla databaser som du har registrerat i %PRODUCTNAME.  
Definiera  
Med den här kommandoknappen definierar du tilldelningen av den nya databasen.  
Så byter du ut en databas i ett dokument mot en annan  
Fältnamn och fälttyper måste vara lika i de båda databaserna om fältkommandona för infogning av datafält ska ge önskade resultat även efter bytet.  
Öppna det dokument där du vill byta ut databasfältkommandon.  
Öppna t.ex. ett nytt dokument baserat på mallen "Affärsbrev", enligt beskrivningen under Skapa standardbrev (kopplad utskrift).  
Öppna dialogrutan Byt databas med kommandot Redigera - Byt databas....  
I vänster listruta, Använda databaser, markerar Du den databastabell som Du vill ersätta och som alltså kommer att skrivas över.  
I höger listruta, Tillgängliga databaser, markerar Du den tabell som ska införas i dokumentet och vars innehåll ska ersätta det hittillsvarande innehållet.  
Klicka på Definiera.  
Du kan kontrollera resultatet av åtgärden med menykommandot Visa - Fältkommandon.  
Infoga (fil)  
Med den här funktionen infogar du en textfil vid markörens position.  
När du har startat den här funktionen visas en dialogruta där du väljer en fil, precis som i dialogrutan Öppna.  
När du har valt en fil, infogas filens innehåll vid markörens position i det aktuella dokumentet.  
Infoga skript  
Med den här funktionen infogar du ett skript vid markörens position i ett text - eller HTML-dokument.  
Om du redan har infogat och markerat ett skript, heter den här dialogrutan Redigera skript.  
Det infogade skriptet indikeras med en liten grön kvadrat i textområdet om du har markerat under Verktyg - Alternativ - HTML-dokument - Vy att anteckningar ska visas.  
Om du dubbelklickar på den lilla gröna kvadraten, öppnas dialogrutan Redigera skript.  
I dialogrutan Redigera skript kan du läsa och redigera skriptets aktuella innehåll.  
Utseendet på dialogrutan Redigera skript skiljer sig från dialogrutan Infoga skript genom två kommandoknappar, med vilka Du kan hoppa mellan föregående respektive följande skript i dokumentet.  
Dessa kommandoknappar syns först om Du har infogat minst två skript i dokumentet.  
Om Du vill kan Du inkludera skriptet vid utskrift, antingen nederst på sidan eller sist i dokumentet.  
Den inställningen gör Du under Arkiv - Skriv ut... - Fler....  
Innehåll  
Skripttyp  
Här anger du skripttyp.  
Skripttypen visas enligt mönstret <SCRIPT LANGUAGE=" JavaScript "> i HTML-koden.  
URL  
Om du vill ange ett länkat skript klickar du på URL och anger skript-filens URL eller väljer filen med hjälp av kommandoknappen till höger.  
HTML-syntaxen för detta är:  
<SCRIPT LANGUAGE=" JavaScript "SRC="url ">  
/* allt här ignoreras * /  
< / SCRIPT>  
...  
Om du klickar på den här kommandoknappen öppnas en dialogruta där du kan infoga en URL.  
Text  
Mata in skriptets text.  
Infoga horisontell linje  
Med den här funktionen infogar du en horisontell linje vid markörens position.  
De horisontella linjerna är identiska med de grafikobjekt som finns i Gallery -temat Linjaler.  
Om du lägger till fler filer i temat Linjaler i Gallery visas även dessa i den här dialogrutan.  
Urval  
Här kan Du välja en linjetyp.  
Sedan klickar Du på OK och linjen infogas.  
Sidhuvud  
På undermenyn till det här kommandot väljer du en sidformatmall i det aktuella dokumentet, vilken ska få ett nytt sidhuvud eller vars sidhuvud du vill ta bort.  
Om du har ett helt nytt oredigerat dokument framför dig, är bara formatmallen Standard tillgänglig.  
Andra sidformatmallar visas först när de verkligen finns.  
Du måste alltså först definiera nya mallar, exempelvis med hjälp av Stylist, eller ladda ett dokument som redan innehåller olika sidformatmallar.  
Klicka på namnet på den sidformatmall som ska få ett sidhuvud.  
Namnet bockmarkeras då, och alla de sidor i det aktuella dokumentet som är försedda med denna sidformatmall får ett nytt tomt sidhuvud.  
Markören placeras automatiskt i det första av de just skapade sidhuvudena, så att Du kan skriva in texten direkt.  
Texten visas samtidigt i alla sidhuvuden med denna sidformatmall.  
Om sidformatmallen på undermenyn redan har bockmarkerats, finns det redan ett sidhuvud för denna sidformatmall.  
Om Du klickar på posten på undermenyn, tas sidhuvudet, efter en säkerhetsfråga, bort från alla de sidor som har denna sidformatmall.  
Även sidhuvudenas eventuella innehåll raderas.  
Om det finns flera sidformatmallar i dokumentet, kan Du också välja Alla, om Du vill ge alla sidor ett sidhuvud eller ta bort det från dem.  
Mer information om sidhuvuden hittar du under menykommandot Format - Sida - Sidhuvud.  
Sidfot  
På undermenyn till det här kommandot väljer du en sidformatmall i det aktuella dokumentet, vilken ska få en ny sidfot eller vars sidfot du vill ta bort.  
Om du har ett helt nytt oredigerat dokument framför dig, är bara sidformatmallen Standard tillgänglig.  
Det är först när du har definierat fler formatmallar, t.ex. med hjälp av Stylist, eller laddar ett dokument som redan innehåller olika formatmallar, som det visas fler sidformatmallar i undermenyn.  
Klicka på namnet på den sidformatmall som ska få en sidfot.  
Namnet bockmarkeras då, och alla sidor i det aktuella dokumentet som är försedda med denna sidformatmall får ett ny tom sidfot.  
Markören placeras automatiskt i den första av de just skapade sidfötterna, så att Du kan skriva in texten direkt.  
Texten visas samtidigt i alla sidfötter med denna sidformatmall.  
Om sidformatmallen på undermenyn redan har bockmarkerats, finns det redan en sidfot för denna sidformatmall.  
Om Du klickar på posten på undermenyn, tas sidfoten, efter en säkerhetsfråga, bort på alla sidor som har denna sidformatmall.  
Även sidfötternas eventuella innehåll raderas.  
Om det finns flera sidformatmallar i dokumentet, kan Du också välja Alla, om Du vill ge alla sidor en sidfot eller ta bort sidfoten från dem.  
Mer information om sidfötter hittar du under menykommandot Format - Sida - Sidfot och i Användarhandboken.  
Fältkommando  
Här kan du infoga fältkommandon i dokumentet.  
På undermenyn kan du direkt välja fält som ofta används.  
Om det önskade fältkommandot inte finns med, väljer du Andra och väljer sedan bland alla tillgängliga fältkommandon.  
Andra...  
Textflöde  
Under den här fliken kan du bestämma hur avstavning och styckebrytning ska göras.  
Avstavning  
I det här området ställer du in egenskaperna för avstavningen i %PRODUCTNAME Writer.  
Automatisk  
Det här alternativet aktiverar den automatiska avstavningen för det aktuella stycket respektive de markerade styckena.  
från... tecken i slutet av raden  
Ange hur många tecken av det avstavade ordet som minst måste finnas kvar i slutet av raden före avstavningen.  
från... tecken i början av raden  
Ange hur många tecken av det avstavade ordet som minst måste finnas på den rad som följer efter avstavningen.  
Högsta antal bindestreck efter varandra  
Ange det maximala antalet på varandra följande rader som får avslutas med ett bindestreck.  
Med 0 görs inga avstavningar.  
Tillägg  
I det här området bestämmer du hur ett stycke ska hanteras om en sidbrytning hamnar i själva stycket.  
Med funktionerna efter rutan Brytning anger du om en sid - eller kolumnbrytning ska infogas före eller efter stycket.  
Brytning  
Med den här kryssrutan aktiverar Du styckebrytning.  
Välj typ av brytning med följande alternativfält.  
Sida  
Om du väljer det här alternativfältet infogas en sidbrytning vid styckebrytningen.  
Kolumn  
Om Du väljer det här alternativfältet infogas en kolumnbrytning vid styckebrytningen.  
Före  
Med det här alternativet infogar Du en sid - eller kolumnbrytning före stycket, och stycket hamnar i början av nästa sida eller kolumn.  
Efter  
Med det här alternativet infogar Du en sid - eller kolumnbrytning efter stycket, och nästa stycke hamnar i början av nästa sida eller kolumn.  
Med sidformatmall  
Aktivera den här rutan om en viss sidformatmall eller ett visst sidnummer ska användas efter sidbrytningen.  
Sidformatmall  
Här väljer du sidformatmall.  
Sidnummer  
I det här rotationsfältet anger Du det sidnummer som Du vill att sidnumreringen ska börja med efter den automatiska sidbrytningen.  
Numret noll (0) betyder att sidnumreringen inte ska ändras.  
Dela inte stycke  
Hela stycket förs odelat över till början av nästa sida eller nästa kolumn om den automatiska sid - eller kolumnbrytningen hamnar inuti stycket.  
Håll ihop stycken  
Det aktuella stycket och nästföljande stycke hålls samman på samma sida eller i samma kolumn.  
Änkekontroll  
Här anger Du hur många rader som minst måste finnas kvar längst ned på sidan för att undvika s k änkor.  
Om det värde som Du anger för rader underskrids, placeras stycket helt och hållet i början på nästa sida.  
Horungekontroll  
Här anger Du hur många rader som minst måste hamna överst på sidan för att undvika s k horungar.  
Om det värde som Du anger för rader underskrids, bryts stycket så att angivet antal rader hamnar överst på nästa sida.  
Anfanger  
Här kontrollerar du anfangsfunktionen för stycket.  
Du anger antal tecken, deras höjd, avståndet från texten och vilken formatmall som ska användas.  
Det eller de första tecknen i början av ett stycke förstoras så att de sträcker sig över flera rader.  
Sådana tecken kallas anfanger.  
Du kan också använda egna tecken (t.ex. symboler) som infogas som anfanger i det markerade stycket.  
Inställningar  
I detta område anger Du inställningarna för anfangsfunktionen i tillämpningsprogrammet.  
Visa anfanger  
Med det här alternativet aktiverar du visningen av anfanger.  
Du får tillgång till alla andra inställningsmöjligheter om du markerar rutan Visa anfanger.  
Helt ord  
Den här rutan är kopplad till Visa anfanger och anger att det första ordet i stycket ska visas som anfang.  
Antal tecken  
Här definierar du hur många tecken i det första ordet i stycket som ska utgöra anfang.  
Rader  
Här definierar du över hur många rader anfangen ska sträcka sig.  
Du kan ange mellan två och nio rader.  
Avstånd till text  
Här anger du avståndet mellan radens början och anfangen.  
Innehåll  
Här kan Du ändra anfangstexten och formatet.  
Anfangstext  
Här inför Du de tecken som ska visas som anfangstext i stället för de första tecknen i styckets början.  
Du kan t ex skriva in symboler, om Du som teckenmall väljer en mall med motsvarande symbolteckensnitt.  
Teckenformatmall  
Här väljer Du en befintlig teckenformatmall.  
Om Du väljer Ingen används det aktuella teckensnittet med aktuella attribut.  
Numrering  
Under den här fliken kan du ställa in en numreringsformatmall vid stycket.  
Dessutom kan du definiera att numreringen ska börja om för det aktuella stycket om du öppnar fliken via dialogrutan Stycke.  
Dessutom kan du styra en radnumrering vid stycket här.  
Du kan börja en numrering vid valfria stycken inom ett dokument eller börja om på nytt.  
Du kan alltså lägga in olika numreringar, som alla har samma formatering, i ett dokument.  
Då kan Du också integrera tabeller, så att numreringen görs, startar eller fortsätter i en tabell.  
Om du ändrar en numrering via Stylist, d.v.s. redigerar stycke - eller numreringsformatmallen, påverkar ändringen alla stycken som är formaterade med respektive mall.  
Men om du ändrar numreringen via dialogrutan Stycke eller dialogrutan Numrering / punktuppställning eller med ikonerna på objektlisten vid numreringar, gör du en direkt formatering och ändringen påverkar bara de stycken i dokumentet som denna formatering används på.  
Numreringsformatmall  
Här väljer Du en numreringsformatmall för stycket.  
Dessa mallar listas även i Stylist, om Du där klickar på ikonen Numreringsformatmallar.  
Numrering  
I det här området kan Du börja om med numreringen av styckena genom att skriva in ett nytt värde för numreringen av det aktuella stycket.  
Det här området visas bara när Du redigerar det aktuella styckets egenskaper, t ex via Format - Stycke..., inte när Du redigerar styckeformatmallen.  
Börja om vid detta stycke  
Markera den här rutan, om Du vill börja en ny numrering vid det aktuella stycket.  
Börja med:  
Här anger Du startvärdet för den nya numreringen.  
Alla följande stycken numreras fortlöpande, såvida Du inte skriver in ett nytt startvärde eller ändrar numreringsformatmallen.  
Radnumrering  
I det här området kan Du göra inställningar för en radnumrering.  
Om Du har aktiverat radnumreringen, kan Du här göra en individuell anpassning av stycket till radnumreringen.  
Räkna med raderna i det här stycket  
Om Du markerar den här kryssrutan, tas raderna i det aktuella stycket med vid en radnumrering.  
Om Du avmarkerar den här rutan, tas inte stycket med vid radnumreringen.  
Börja om vid detta stycke  
Om den här kryssrutan är markerad, börjar en radnumrering om vid det aktuella stycket.  
Om Du vill kan Du ange ett startvärde.  
Börja med:  
Här kan Du ange med vilket startvärde en radnumrering ska börja om vid stycket.  
Sidformatmall  
Med den här funktionen kan du definiera utseendet för hela sidan.  
Du bestämmer bl.a. marginaler, pappersformat, stående och liggande format, sidhuvuden och sidfötter, indelning i kolumner och placeringen av fotnoter.  
Dessutom kan du bestämma vilken inramning och bakgrund sidorna ska ha här.  
Kolumner  
Här kan du definiera antalet kolumner per sida, ram eller område.  
Vidare kan du bestämma typ, höjd och placering för linjen mellan kolumnerna samt ändra kolumnbredden.  
Förinställningar  
I detta område anger Du antalet kolumner.  
Dessutom kan Du välja kolumnlayout bland dem som visas i exempelrutorna.  
Kolumninställningarna för sidor gäller alla de sidor där den aktuella sidformatmallen används.  
Kolumninställningarna för flerkolumniga ramar gäller den aktuella ramen eller - vid ändring av ramformatmallen - alla ramar som baseras på den mallen (eller en mall som är baserad på den).  
Kolumner  
Här anger Du antal för de kolumner som ska skapas i textområdet mellan sidomarginalerna eller vänster och höger ramkant.  
Du behöver inte ange ett kolumnantal utan kan välja kolumnlayouten i något av de fem valfälten genom att markera den.  
Urvalsfält  
Här kan du välja bland ofta använda standardinställningar.  
Fördela innehåll jämnt över alla kolumner  
Om den här rutan är markerad, fördelas textinnehållet i områden med flera kolumner så jämnt som möjligt mellan kolumnerna.  
Annars fylls kolumnerna löpande ut med text från den första till den sista kolumnen.  
Bredd och avstånd  
Du kan bara ändra kolumnbredd om rutan Automatisk bredd inte är markerad.  
(Kolumnnummer)  
Här visas kolumnnumren.  
Därunder står kolumnbredden och avståndet till intilliggande kolumner.  
Vänsterpil  
Vid fler än tre kolumner kan Du visa de kolumner som står till vänster om visningsområdet med hjälp av den här symbolen.  
Vänsterpil  
Högerpil  
Vid fler än tre kolumner kan Du visa de kolumner som står till höger om visningsområdet med hjälp av den här symbolen.  
Högerpil  
Bredd  
I rotationsfälten kan du ändra bredden på kolumnen vars nummer visas ovanför fältet.  
Du kan bara använda rotationsfälten om rutan Automatisk bredd inte är markerad.  
Avstånd  
Här definierar du avståndet mellan de båda kolumnerna som visas ovanför.  
Automatisk bredd  
Om du vill att kolumnerna ska ha samma bredd, markerar du den här rutan.  
Vid förhandsgranskningen av en flerkolumnig textram visas bara kolumnindelningen inom ramen, inte den omgivande sidan.  
Skiljelinje  
Det här området är aktivt bara om antalet kolumner är minst två.  
Du kan skilja kolumnerna åt med skiljelinjer.  
Typ  
Här kan Du välja mellan olika linjebredder.  
Om Du inte vill ha någon skiljelinje mellan kolumnerna väljer Du Ingen.  
Höjd  
Du kan bara använda det här rotationsfältet om Du har valt en linjebredd i fältet Typ.  
Här anger Du skiljelinjens höjd i förhållande till textområdets höjd.  
Som standard anges en skiljelinje som går från topp - till bottenmarginal.  
Position  
Listrutan är tillgängligt bara om värdet i fältet Höjd är mindre än 100%.  
Du kan välja mellan positionerna Överst, Centrerad och Nederst.  
Använd på  
När du har valt kommandot Format - Kolumner, väljer du här om redigeringen av kolumnerna ska tillämpas på det valda textavsnittet (d.v.s. där markören står) eller på sidformatmallen.  
Alternativ  
Här kan Du definiera antalet textkolumner och bakgrunden i det infogade området.  
Du kan också bestämma typ, höjd och placering av kolumnernas skiljelinje och ändra kolumnbredden.  
Områden i StarWriter kan nu innehålla kolumner.  
Områdena underordnar sig textflödet på den plats i dokumentet, där de har infogats.  
Det innebär för det första att om Du infogar ett område med kolumner på en sida, vilken i sin tur är uppdelad i kolumner, får Du kolumner inuti kolumnerna.  
Områdets kolumner ligger innanför sidans kolumner.  
För det andra kan Du infoga ett område i ett annat område.  
Om båda områdena har kolumner, avbryts bara det överordnade områdets kolumnuppdelning och fortsätter när det underordnade området har upphört.  
Möjligheten att kunna definiera kolumner i områden gör det lättare att importera och exportera till andra program, där flera olika kolumnuppdelningar per sida är möjliga.  
För närvarande stöds denna funktion vid import och export i RTF-format, import i Word-format och import i WordPerfect8-format.  
Även export i Word-format kommer inom kort att utökas med denna funktion.  
Fotnot  
Under fliken Fotnot definierar du var på sidan fotnoter är tillåtna och typen av skiljelinje.  
Om den här fliken inte visas, har Du aktiverat läget Utskriftslayout.  
Då visas inte fotnoter.  
Fotnotsområde  
Här definierar Du fotnotsområdets höjd.  
Höjd maximalt som sidan  
Markera det här alternativfältet om Du vill att höjden på fotnotsområdet automatiskt ska anpassas efter antalet fotnoter.  
Fotnotens max höjd  
Om Du vill begränsa storleken på fotnotsområdet klickar Du här.  
Fotnotens max höjd  
Det här rotationsfältet kan Du enbart använda om Du har markerat alternativfältet Fotnotens max höjd.  
Här anger Du maximal höjd på fotnotsområdet.  
Avstånd från brödtext  
Här anger Du avståndet mellan bottenmarginalen och första textraden i fotnotsområdet.  
Löptexten förskjuts uppåt i motsvarande mån.  
Skiljelinje  
I det här området väljer Du skiljelinjens placering och längd.  
Position  
Här anger Du den horisontella justeringen av skiljelinjen mellan fotnotsområdet och brödtexten.  
Längd  
I det här rotationsfältet anger Du över hur många procent av textområdet skiljelinjen ska sträcka sig.  
Styrka  
Här väljer Du önskad linjebredd på skiljelinjen.  
Avstånd till fotnotens innehåll  
Här anger Du avståndet mellan fotnotsområdet och skiljelinjen.  
Löptexten förskjuts uppåt i motsvarande mån.  
Avståndet mellan två fotnoter ställer Du in under Format - Stycke - Indrag och avstånd.  
I området Avstånd kan Du enkelt ange hur stort avståndet ska vara före respektive efter ett stycke.  
Fot - / slutnoter  
Under fliken Fot - / slutnoter bestämmer du om fotnoter och / eller slutnoter ska samlas vid textslutet och få en egen nummersekvens.  
Om den här fliken inte visas, har du aktiverat utskriftslayouten.  
I det läget är fotnoter inte inlagda.  
Fotnoter  
Definiera här var fotnoter placeras i områden.  
samla vid textslut  
Markera den här rutan, om fotnotens innehåll ska placeras i slutet av området eller i slutet av sidan.  
Fotnoten placeras i slutet av sidan om området fortsätter på följande sida.  
oberoende numrering  
Om du vill infoga en egen numrering för fotnoterna, markerar du den här rutan.  
Börja med  
Välj här med vilket nummer numreringen ska börja.  
eget format  
Om du vill använda en annan numrering än den som angetts under oberoende numrering / Börja med, klickar du i den här rutan.  
Den är bara tillgänglig om rutan oberoende numrering har markerats först.  
Före  
Tecknen som har skrivits in i det här textfältet placeras framför numreringen.  
Rotationsfält eget format  
Här väljer du lämplig numrering för fotnoterna.  
Efter  
I textfältet kan du skriva in tecken som ska infogas efter fotnotsnumreringen.  
Slutnoter  
Här definierar du var slutnoter ska placeras i områden.  
samla vid områdets slut  
Markera den här rutan, om slutnotens innehåll ska placeras vid områdets slut.  
oberoende numrering  
Om du vill infoga en egen numrering för slutnoterna, markerar du den här rutan.  
Börja med  
Välj här med vilket nummer slutnotsnumreringen ska börja.  
eget format  
Om du vill använda en annan numrering för slutnoterna än den som är förinställd under oberoende numrering / Börja med, markerar du den här rutan.  
Den är bara tillgänglig om rutan oberoende numrering har markerats först.  
Före  
Tecknen som du skriver in i det här textfältet placeras före slutnotsnumreringen.  
Rotationsfält eget format  
Här väljer du lämplig numrering för slutnoterna.  
Efter  
I textfältet kan du skriva in tecken, som ska infogas efter slutnotsnumreringen.  
Grafik  
Med den här funktionen redigerar du egenskaperna för ett grafikobjekt.  
Du kan också redigera ett markerat grafikobjekt med särskilda kortkommandon.  
Dialogrutan Grafik öppnas med följande flikar:  
Textanpassning  
Typ  
Under den här fliken definierar du storlek och placering för ett objekt på sidan.  
Det kan vara en ram, ett grafikobjekt eller ett annat objekt.  
Storlek  
Här bestämmer du storleken på objektet.  
Bredd  
I det här rotationsfältet anger Du objektets bredd.  
Relativ  
Om Du markerar det här alternativet, kan Du i rotationsfältet Bredd ange objektets relativa bredd.  
I online-layouten hänför sig den relativa bredden till sidbredden, i tabellceller till cellens bredd, och i en ram är den bredden på ramens utskriftsområde.  
I alla andra fall används sidans utskriftsområde som relativ referens.  
Höjd  
Här kan Du ändra objektets höjd.  
Relativ  
Om Du markerar det här alternativet, kan Du ange objektets höjd i förhållande till höjden på sidans utskriftsområde i rotationsfältet Höjd.  
Anpassa proportionellt  
Om Du markerar den här kryssrutan, blir varje förändring av objektet proportionell.  
Detta kan vara nödvändigt för att t ex undvika att bilder förvrids.  
Originalstorlek  
Klicka här om Du vill upphäva storleksändringar och återgå till objektets originalstorlek.  
Om Du redigerar en ram, visas inte den här kommandoknappen.  
Automatisk höjd  
Markera den här kryssrutan när Du vill att ramens höjd automatiskt ska anpassas till den text som den innehåller.  
Om kryssrutan inte är markerad och texten sträcker sig längre än ramens underkant, kommer texten nedanför kanten inte att synas.  
Den här kryssrutan visas bara när Du redigerar en ram.  
Förankring  
Välj typ av förankring för objektet här.  
Mer information hittar Du under Format - Förankring.  
Vid sidan  
Med det här alternativet kopplar du objektet till den aktuella sidan.  
Vid stycke  
Med det här alternativet kopplar du objektet till det aktuella stycket.  
Vid tecken  
Med det här alternativet kopplar du objektet till ett tecken.  
Som tecken  
Med det här alternativet uppför sig objektet som ett tecken: det står som en vanlig bokstav i textflödet och påverkar radhöjd och radbrytning på samma sätt som en bokstav.  
Eftersom objektets horisontella position bestäms av textflödet, kan du under Position bara ställa in den vertikala justeringen med avseende på den aktuella raden.  
Position  
I det här området kan Du ändra objektets placering.  
Placeringsangivelsen är alltid relativ, varvid de olika referenselementen kan vara t ex marginaler eller styckekanter, och den beror på förankringens typ.  
Mer information hittar Du under Format -Justering.  
Horisontellt  
Här anger Du alternativet för den horisontella justeringen.  
I kombinationsfältet till anger Du det referenselement som justeringen ställs in efter.  
Denna funktion är inte tillgänglig för Förankring som tecken.  
med  
Här anger Du det horisontella avståndet mellan vänster kant på det referenselement som Du har valt i kombinationsfältet till och vänster kant på det objekt som ska justeras.  
Rotationsfältet är aktivt bara om Du har valt alternativet Från vänster i kombinationsfältet Horisontellt.  
till  
Här anger Du det referenselement som objektets horisontella justering ska hänföra sig till.  
De olika alternativen beror på förankringens typ.  
Vid förankring till sidan, till ett stycke och till ett tecken kan Du göra en horisontell justering i förhållande till sidmarginalerna, hela sidan eller sidtextområdet.  
När Du förankrar till ramen kan Du på motsvarande sätt göra justeringen i förhållande till en ramkant, hela ramen eller ramtextområdet.  
För ramar som är kopplade till stycke och förankrade till tecken finns det ytterligare referenselement, nämligen styckemarginaler, styckeområde och textområde i stycke.  
Textområdet på sidan motsvarar i allmänhet styckeområdet; dock gäller inte detta sidor med flera kolumner.  
Textområdet i stycke är stycke( området) utan styckekanter; på motsvarande sätt är textområdet på sidan själva sidan utan sidmarginaler och ramtextområdet i ramen utan ramkanter.  
De olika definitionerna visas om Du väljer respektive referenselement i förhandsvisningsfältet.  
spegelvänt på jämna sidor  
Om den här kryssrutan är aktiv, spegelvänds inställningarna för den horisontella justeringen på jämna sidor.  
Det innebär att justeringsoperationerna Vänster, Höger eller Från vänster utvärderas spegelvänt på jämna sidor.  
Om Du exempelvis justerar objektet vänsterställt på en udda sida, kommer det att efter en sidbrytning justeras högerställt på nästa sida.  
Justeringsalternativen heter därför Invändigt i stället för Vänster och Utsida i stället för Höger.  
Speglingen gäller både objektets justering och för referenselementet.  
På detta sätt kan Du skapa exempelvis en ram eller ett grafiskt objekt som alltid befinner sig i innerkanten på sidans yttermarginal.  
Om det är ett grafikobjekt som ska justeras, t ex en pil, kan Du dessutom använda speglingsalternativet Sidor, om Du inte bara vill anpassa objektets placering utan även hur dess innehåll ska visas på udda och jämna sidor.  
Vertikalt  
Här anger Du alternativet för den vertikala justeringen.  
I kombinationsfältet till anger Du det referenselement som justeringen ställs in efter.  
När du förankrar vid en ram bör du lägga märke till att alternativen Nederst och Mitten bara är tillgängliga för vertikal justering om den omgivande ramen har fast höjd.  
Om höjden på den omgivande ankarramen automatiskt anpassas till sitt innehåll (kryssrutan Automatisk höjd), kan du bara justera den infogade ramen mot överkanten på den omgivande ramen.  
med  
Här anger Du det vertikala avståndet mellan det referenselement som Du har valt i kombinationsfältet till och överkanten på det objekt som ska justeras.  
Det här rotationsfältet är aktivt bara om Du i kombinationsfältet Vertikalt har valt alternativet Uppifrån eller, vid förankring som tecken, Nedifrån.  
Vid alternativet Uppifrån anger Du avståndet till överkanten på referenselementet; vid alternativet Nedifrån och förankring som tecken anger Du avståndet till baslinjen.  
till  
Här anger Du det referenselement som objektets vertikala justering ska hänföra sig till.  
De olika alternativen beror på förankringens typ.  
Om Du har valt Förankring som tecken, kan Du välja mellan referenselementen Baslinje, Tecken och Rad.  
Vilka effekter de olika alternativen har visas i förhandsvisningsfältet.  
I förhandsvisningen visas den som en röd linje.  
Alternativet Tecken står för den höjd som alla tecken på raden (inklusive staplar) har.  
Alternativet Rad står för den fullständiga radhöjden inklusive alla objekt som är kopplade som tecken.  
Ett tvådimensionellt referenselement som justeringen hänför sig till visas som en röd kvadrat och det justerade objektet som en grön.  
Baslinjen utmärks med en röd linje om objektet förankras som tecken.  
Textanpassning  
Här kan du definiera textanpassningen kring ett objekt.  
Det kan t.ex. vara en ram, ett grafikobjekt eller en teckning.  
Vidare kan du definiera objektets placering vid sidväxling samt avstånden mellan text och objekt.  
Om du vill ha textanpassning runt en texttabell sätter du texttabellen i en ram och definierar sedan textanpassningen runt ramen.  
Förinställningar  
I det här området definierar du hur text och objekt ska förhålla sig till varandra.  
Ingen  
Välj det här alternativet när texten ska avbrytas av ramen, det grafiska objektet eller objektet.  
Texten slutar då ovanför objektet, oavsett hur brett objektet är, och fortsätter sedan nedanför det.  
Det är tomt på båda sidor om objektet.  
Ingen  
Vänster  
Om det finns fritt utrymme till vänster om objektet löper texten där.  
Vänster  
Höger  
Om det finns fritt utrymme till höger om objektet löper texten där.  
Höger  
Parallell  
Texten löper till vänster och höger om objektet om det finns tillräckligt med plats.  
Varje rad avbryts då av objektet.  
Parallell  
Genomflöde  
Välj det här alternativet när texten ska flöda bakom ramen, det grafiska objektet eller objektet.  
Objektets innehåll täcker då texten.  
Genomflöde  
Dynamisk  
Texten löper runt objektet till höger, vänster eller inte alls beroende på det utrymme som finns.  
Om avståndet mellan objekt och marginal är mindre än 2 cm, hamnar dock ingen text där.  
För objekt vars bredd underskrider 1,5 cm och där avståndet till marginalerna är större än 2 cm, blir textanpassningen parallell.  
Dynamisk  
Alternativ  
Här anger Du alternativen för textanpassning.  
Första stycket  
Aktivera den här funktionen när du har tryckt på Retur och sedan vill påbörja ett nytt stycke nedanför objektet.  
Avståndet mellan styckena avgörs av objektets storlek.  
Med det här alternativet kan du t.ex. se till att det aktuella stycket, vid vilket objektet är förankrat, löper runt om objektet medan det följande stycket, som kanske är en rubrik, inte placeras bredvid objektet utan nedanför det.  
I bakgrunden  
Objekt och text överlappar varandra.  
Det här alternativet är bara tillgängligt om du har valt textanpassningstypen Genomflöde.  
Kontur  
Om du väljer den här funktionen, flyter texten runt objektets kontur.  
Funktionen är särskilt effektfull för polygoner.  
Om du har valt textanpassningen Genomflöde kan du inte välja den här funktionen. %PRODUCTNAME känner igen de flesta konturer automatiskt.  
I Konturredigeraren kan du anpassa konturen som du vill manuellt.  
Konturredigeraren öppnar du genom att välja menykommandot Textanpassning på formatmenyn till ett infogat grafikobjekt, och därefter menykommandot Redigera kontur Du kan också välja det här menykommandot på snabbmenyn till ett infogat grafikobjekt.  
Infogade 3D-objekt kan du också förse med konturanpassningar.  
Genom att kombinera detta med att låta text flyta inuti objekt, kan du åstadkomma imponerande effekter.  
Objekt som du ändrar på detta sätt kan du förstås även lägga in i presentationer.  
Den här funktionen är inte tillgänglig för ramar.  
Bara utanför  
När Du har valt konturanpassning, kan Du med det här alternativet ange att texten bara ska flöda till vänster och höger om objektet men inte "inuti".  
Texten avbryts alltså högst en gång av objektet.  
Det här alternativet kan Du inte använda för ramar.  
Avstånd  
I det här området anger Du de enskilda avstånden mellan objektets kant och texten.  
Avstånden gäller mellan texten och objektets ytterkant när Du har aktiverat konturanpassningen mellan texten och objektets kontur i angiven riktning.  
Lägg märke till att Du kan ange avstånden till vänster, höger, ovanför och nedanför var för sig, och att de också hänför sig till text som löper inuti objektet, såvida Du inte har ställt av konturanpassning inuti objektet.  
Skriv t ex versala initialer i %PRODUCTNAME Impress, omvandla dem till kurvor, kopiera dem till Urklipp och infoga dem i ett textdokument.  
Vänster  
Här definierar Du avståndet mellan objektets vänsterkant och texten.  
Höger  
Här definierar Du avståndet mellan objektets högerkant och texten.  
Överst  
Här definierar Du avståndet mellan objektets övre kant och texten.  
Underst  
Här definierar Du avståndet mellan objektets nedre kant och texten.  
Konturredigerare  
Här redigerar du konturerna för grafik, objekt och ramar.  
Dessa konturer gäller för kontur-textanpassningen.  
I visningsfältet visas det redigerade grafikobjektet och de konturer som Du har definierat.  
Tilldela  
Efter varje ändring i konturredigeraren klickar du på den här ikonen för att tilldela den aktuella ändringen.  
Tilldela  
Arbetsområde  
Klicka här om du vill radera den befintliga konturen och definiera ett nytt arbetsområde.  
Arbetsområde  
Urval  
Klicka på symbolen Urval så aktiveras urvalsmarkören.  
Med den här markören kan Du klicka på en annan del i konturen för att sedan redigera den.  
Urval  
Rektangel  
Klicka på Rektangel om Du vill definiera ett rektangulärt område.  
Markören får en liten rektangel bredvid hårkorset och Du kan nu dra ut en rektangel.  
Om Du vill skapa en kvadrat håller Du ned skifttangenten samtidigt som Du drar.  
Rektangel  
Ellips  
Klicka på Ellips om Du vill definiera ett runt område.  
Markören får en liten cirkel bredvid hårkorset och Du kan nu dra ut en ellips.  
Om Du vill skapa en cirkel håller Du ned skifttangenten samtidigt som Du drar.  
Ellips  
Polygon  
Klicka på Polygon om Du vill definiera ett valfritt område.  
Markören får en liten kurva bredvid hårkorset och Du kan nu definiera en polygon.  
Klicka på varje punkt på kurvan som Du vill definiera.  
Dubbelklicka på startpunkten för att sluta kurvan.  
Du kan begränsa vinkeln till multipler av 45 grader om Du håller ned skifttangenten när Du placerar muspekaren.  
Polygon  
Redigera punkter  
Klicka på Redigera punkter om Du vill visa enstaka stödpunkter på Bézierkurvor.  
Då kan Du redigera de enskilda stödpunkterna på kurvan med hjälp av musen.  
Redigera punkter  
Flytta punkter  
Klicka på Flytta punkter om Du vill flytta enstaka punkter som definierar en polygon.  
Flytta punkter  
Infoga punkter  
Klicka på Infoga punkter om Du vill infoga ytterligare stödpunkter.  
Infoga punkter  
Radera punkter  
Klicka på Radera punkter om Du vill ta bort enstaka stödpunkter.  
Radera punkter  
AutoKontur  
Om Du klickar på den här ikonen skapar Du en kontur runt objektet som Du sedan kan finjustera.  
AutoKontur  
Ångra  
Med den här kommandoknappen ångrar Du den senast utförda åtgärden.  
Ångra  
Upprepa  
Med den här kommandoknappen upprepar Du den senast utförda åtgärden.  
Upprepa  
Pipett  
Här aktiverar Du pipetten för bitmapbilder.  
Klicka på en färg på bitmapbilden med pipetten.  
Alla pixlar som är direkt förbundna med pixeln som Du har klickat på och som har samma färg sammanfattas till en kontur.  
Som "samma" färg räknas de färger som ligger inom det toleransområde som Du ställer in med rotationsknapparna.  
Vid 0% tolerans måste färgen stämma exakt överens och med 100% tolerans gäller alla färger som samma färg.  
Pipett  
Färgtolerans  
I det här rotationsfältet kan Du ställa in den önskade färgtoleransen för pipetten.  
Grafik  
Här kan du spegelvända ditt grafikobjekt samt uppdatera länken till en grafikfil.  
Spegelvänd  
I det här området kan du spegelvända grafikobjektet horisontellt och vertikalt.  
Mer information finns under Format - Spegelvänd.  
vertikalt  
Med det här alternativet spegelvänder du grafikobjekt vertikalt.  
Det kan du också göra med ikonen på objektlisten.  
horisontalt, på  
Med det här alternativet spegelvänder du grafikobjektet horisontellt.  
I det tillhörande alternativfältet väljer du om ett grafikobjekt ska spegelvändas likadant på alla sidor eller bara på höger - resp. vänstersidor.  
Du kan även använda ikonen på objektlisten.  
på alla sidor  
När du spegelvänder horisontellt kan du här välja om grafikobjektet ska vara spegelvänt horisontellt på alla sidor, eller bara på vänster - eller på högersidor.  
på vänstersidor  
Här kan du välja om grafikobjektet ska spegelvändas horisontellt på vänstersidor.  
på högersidor  
Här kan du välja om grafikobjektet ska spegelvändas horisontellt på högersidor.  
Länk  
I det här området kan du uppdatera länkningen till en grafikfil.  
Mer information finns under Redigera - Länkar.  
Filnamn  
Om grafikobjektet är infogat som länk, står den fullständiga sökvägen till den länkade filen här.  
Du kan ändra sökvägen direkt med tangenterna eller genom att klicka på kommandoknappen....  
...  
Med den här kommandoknappen öppnar du dialogrutan Länka.  
Där kan du välja en annan grafikfil eller uppdatera sökvägen till den önskade grafikfilen.  
Dialogrutan Länka är uppbyggd på samma sätt som dialogrutan Infoga grafik.  
Makro  
Här kan du välja ett makro som ska utföras vid en viss händelse.  
Därmed är händelsen kopplad till det aktuella objektet.  
Beroende på objektet hittar du den här funktionen under fliken Makro i respektive objektdialogruta eller i dialogrutan Tilldela makro.  
Händelse  
Här listas händelserna tillsammans med de aktuella tilldelade makrokommandona.  
Bara de alternativ som är definierade för det aktuella objektet visas.  
För alla objekt som är infogade i ett dokument och som kan kopplas till ett makro visas i den följande tabellen respektive definierade händelser.  
Händelse  
Händelsen inträffar...  
OLE-objekt  
Grafik  
Ram  
AutoText  
ImageMap-area  
Hyperlänk  
Klicka på objekt  
...om objektet markeras.  
x  
x  
x  
Mus över objekt  
... när muspekaren förs över objektet.  
x  
x  
x  
x  
x  
Utför hyperlänk  
... när en hyperlänk-URL har definierats för objektet och hyperlänken aktiveras.  
x  
x  
x  
x  
Mus lämnar objekt  
... när muspekaren förs bort från objektet.  
x  
x  
x  
x  
x  
Laddning av grafik lyckades  
... när grafikobjektet har laddats utan problem.  
x  
Laddning av grafik avbröts  
... när laddningen av grafikobjektet avbröts av användaren (t.ex. vid en nedladdning).  
x  
Fel vid laddning av grafik  
... när laddningen av grafikobjektet inte kunde genomföras (t.ex. därför att det inte kunde hittas).  
x  
Inmatning av alfatecken  
... när inmatning av bokstäver, siffror och andra tecken som textinmatning görs via tangentbordet.  
x  
Inmatning av icke-alfatecken  
... när användaren matar in kontrolltecken från tangentbordet såsom tabbar, radbrytning mm.  
x  
Ändra ramstorlek  
... när användaren ändrar ramens storlek med musen.  
x  
Flytta ram  
... när ramen flyttas med musen.  
x  
Innan AutoText infogas  
... innan ett textblock infogas.  
x  
När AutoText har infogats  
... när ett textblock har infogats.  
x  
Händelser som är bundna till kontrollfält i ett formulär beskrivs i hjälpen till Kontrollfältegenskaper.  
Dem hittar Du i Formuläregenskaperna.  
Makron  
I det här området väljer Du det makro som ska exekveras när en viss händelse inträffar.  
När det gäller ramar kan du koppla vissa händelser till en FUNCTION där du kan bestämma om händelsen ska bearbetas av %PRODUCTNAME Writer eller av denna FUNCTION.  
Mer information finns i %PRODUCTNAME Basic-hjälpen.  
Kategori  
Här förtecknas programmet %PRODUCTNAME och de öppna dokumenten.  
Välj i listan var makrona ska sparas.  
Makronamn  
Här visas namnen på de makron som är tillgängliga på den valda enheten.  
Markera önskat makro.  
Tilldela  
Med hjälp av den här knappen tilldelar Du det makro som Du har markerat i området Makron den händelse som Du har valt under Händelse.  
Uppgifterna om det tilldelade makrot visas efter händelseposten.  
Upphäv  
Med den här kommandoknappen upphäver du tilldelningen av ett makro till den markerade posten i området.  
Du blir inte ombedd att bekräfta åtgärden.  
Urvalsfältet Makron  
I den här listrutan kan du välja att du vill tilldela ett %PRODUCTNAME Basic-makro.  
%PRODUCTNAME Basic  
Klicka på det här alternativet om du vill tilldela ett %PRODUCTNAME Basic-makro.  
Hyperlänk  
Här väljer du hyperlänkegenskaper för grafikobjekt, ramar eller OLE-objekt.  
Länk till  
I det här området anger du den URL som du ska gå till när du klickar på grafikobjektet, objektet eller ramen.  
URL  
Ange här hela URL:en.  
Här följer några exempel: http: / /www.sun.de eller file: / //c _BAR_ / Office / Document / Internet.sdw.  
Välj ut...  
Med den här kommandoknappen öppnar Du dialogrutan Öppna.  
Namn  
Namnge hyperlänkgrafiken i det här fältet.  
Ram  
I det här fältet anger du den målram, där den laddade URL:en ska visas.  
De förinställda posternas betydelse hittar Du i förklaringstabellen.  
Image map  
Här markerar du typen av Image map, som tilldelats grafikobjektet, OLE-objektet eller ramen.  
Inställningarna för URL och målram i området Hyperlänk gäller bara, om du inte skapar någon image map.  
Annars gäller inställningarna för image map.  
Image map på serversidan  
Markera det här alternativet om objektet är en image map på serversidan.  
Image map på klientsidan  
Det här alternativet är markerat, om objektet tilldelats en image map på klientsidan.  
Då måste en Image map ha definierats för detta objekt.  
Tillägg  
Här kan du bestämma och redigera fler egenskaper för en ram, ett grafikobjekt eller ett objekt.  
Namn  
Här kan du redigera namnet på objektet eller bestämma om det ska anges en alternativtext för namnet på ramen, grafikobjektet eller objektet.  
Namn  
I det här området kan du tilldela ramen, grafikobjektet eller objektet ett namn.  
Skriv in ett namn eller använd helt enkelt den föreslagna beteckningen.  
Med hjälp av namnen kan du lättare skilja dem åt.  
De namn som du väljer här visas t.ex. i Navigator.  
När du redigerar långa dokument underlättar det arbetet betydligt om du har tilldelat namn enligt en enhetlig princip.  
Alternativtext (för grafikobjekt och objekt)  
Om du skriver in en text här, visas den om du pekar på ett grafikområde med musen.  
Den här funktionen är bara relevant om du skapar webbdokument.  
Det här textfältet visas bara vid grafikobjekt eller OLE-objekt, inte vid ramar.  
Föregående  
I det här fältet visas namnet på föregående ram, om den är länkad till den aktuella.  
Följande  
I det här fältet visas namnet på efterföljande ram, om den är länkad till den aktuella.  
Skydda  
I det här området kan du ange om och hur ramen i dokumentet ska skyddas mot en ändring.  
Skydda innehåll  
Om du aktiverar den här rutan, skyddas innehållet i ramen och kan inte längre ändras.  
Om markören står i en skrivskyddad ram, visas "skrivskyddad" på statuslisten.  
Du kan t.ex. kopiera raminnehållet men inte klippa ut det.  
Skydda position  
Om du aktiverar den här rutan, kan du inte ändra objektets placering av misstag.  
Skydda storlek  
Om du aktiverar den här rutan kan du inte ändra objektets storlek av misstag.  
Egenskaper  
I det här området hittar du alternativ för att skydda grafikobjekt, ramar eller objekt mot oavsiktliga ändringar.  
Redigerbar i skrivskyddat dokument (bara vid ramar)  
Om du aktiverar den här rutan, kan du redigera innehållet i en ram även om dokumentet är skrivskyddat.  
Skriv ut  
Om du har aktiverat den här rutan, skrivs grafikobjektet, ramen eller objektet också ut.  
Med det här kommandot öppnar du dialogrutan Objekt.  
Här kan du ändra objektets egenskaper, t.ex. storlek, namn, placering, textanpassning, inramning med mera.  
Du kan också ändra ett markerat objekt med särskilda kortkommandon.  
Textanpassning  
Tabellformat  
Med den här funktionen kan du definiera tabellegenskaper.  
Bestäm egenskaper som namn, justering, avstånd, kolumnantal, kolumnbredd, inramning och bakgrund.  
Tabell  
Här kan du definiera tabellens storlek och justering.  
Dessutom kan du definiera avståndet till styckena som omger tabellen.  
Egenskaper  
I det här området kan du definiera tabellegenskaper, t.ex. namn och bredd.  
Namn  
Här anger Du vilket namn tabellen ska ha internt.  
Bredd  
Ange här önskad totalbredd på tabellen.  
Det här rotationsfältet kan Du inte använda om Du har markerat alternativfältet Automatisk.  
Relativ  
Om Du markerar den här kryssrutan, visas tabellbredden i procent av sidbredden.  
Justering  
I det här området anger Du tabellens justering i förhållande till dokumentsidan.  
Automatiskt  
Klicka här om tabellen ska sträcka sig från vänster till höger marginal.  
Detta är den rekommenderade inställningen för tabeller på HTML-sidor.  
Vänster  
Om Du klickar här, placeras tabellen intill vänstermarginalen.  
Du kan själv ange bredden.  
Från vänster  
Om Du vill ställa in ett avstånd från vänstermarginalen och kunna ge tabellen en viss bredd, måste Du först markera det här alternativfältet.  
I fälten Till vänster och Bredd anger Du sedan önskade värden.  
Höger  
Om Du klickar här, placeras tabellen intill högermarginalen.  
Du kan själv ange bredden.  
Centrerat  
Om Du klickar här, placeras tabellen mitt emellan vänster - och högermarginalen.  
Ange tabellens totalbredd eller ange avståndet mellan vänstermarginalen och den första tabellkolumnen i fältet Till vänster.  
Manuellt  
Om Du klickar här, placeras tabellen i enlighet med de gällande värdena i rotationsfälten Till vänster och Till höger mellan vänster och höger marginal.  
Tabellbredden räknas ut automatiskt.  
Det är bara med den här inställningen som Du kan reglera kolumnbredderna oberoende av varandra.  
Avstånd  
I det här området anger Du avstånden till vänster - och högermarginalen och till föregående och efterföljande textstycke.  
Till vänster  
Här anger Du avstånd från vänster marginal till den första tabellkolumnen.  
Den här rotationsrutan kan användas bara om Du har valt något av alternativen Från vänster, Höger eller Manuellt under Justering.  
Till höger  
Här anger Du avståndet från den sista tabellkolumnen till högermarginalen.  
Den här rotationsrutan kan Du bara använda om Du har valt något av alternativen Vänster och Manuellt under Justering.  
Upp  
Här anger Du avståndet mellan den sista raden i textstycket ovanför tabellen och den första raden i tabellen.  
Ner  
Här anger Du avståndet mellan den sista raden i tabellen och den första raden i textstycket nedanför tabellen.  
Om tabellen står först i dokumentet eller i ett sidhuvud eller en sidfot, kan Du infoga ett stycke ovanför tabellen genom att trycka på returtangenten när markören står i den första cellen.  
Om Du vill ta bort ett tomt stycke ovanför en tabell, trycker Du på backstegstangenten när markören står i den första cellen.  
Kolumner  
Här kan du ändra kolumnbredden för alla kolumner i tabellen manuellt.  
Hur du ändrar kolumnbredden med hjälp av mus och tangentbord, utan att behöva öppna en dialogruta, får du reda på under den här hyperlänken:  
Anpassa tabellbredd  
Om den här rutan är markerad, kan alla kolumnbredder i tabellen ändras oberoende av de andra.  
Den här rutan är bara aktiv, om Du har markerat justeringen Manuellt på fliken Tabell.  
Ändra kolumner proportionellt  
Markera den här rutan, om Du vill ändra alla kolumner lika mycket.  
De olika kolumnernas relativa andelar av hela tabellbredden förblir de samma.  
Den här rutan är bara aktiv, om Du har markerat justeringen Manuellt på fliken Tabell.  
Återstående plats  
I det här visningsfältet visas hur mycket plats som finns kvar att tilldela de olika kolumnbredderna tills du har uppnått den totala bredd som du kan ställa in under fliken Tabell.  
Kolumnbredd  
I det här området visas den aktuella kolumnbredden som du kan ändra.  
Om en tabell innehåller mer än sex kolumner, kan du växla till de kolumner som inte visas med hjälp av pilknapparna.  
Kolumnbredder  
I dessa rotationsfält definierar Du den nya kolumnbredden.  
Om Du ändrar en kolumnbredd inverkar det nästan alltid på bredden på nästa kolumn.  
Ändringar av den sista kolumnen inverkar på den första tabellkolumnen.  
Detta gäller inte om Du har markerat kryssrutan Anpassa tabellbredd.  
Då kan Du ändra varje kolumn oberoende av de övriga.  
Vänsterpil  
Om tabellen skulle innehålla fler än sex kolumner, kan Du här växla till de kolumner till vänster som inte visas.  
Högerpil  
Här kan Du växla till de kolumner till höger som inte visas.  
Redigera tabell via tangentbord  
Här följer en kort beskrivning av hur du kan redigera en tabell i ett textdokument med hjälp av tangentbordet.  
Flertalet av de funktioner som beskrivs här kan du även nå via objektlisten för tabeller eller snabbmenyn.  
Flytta kolumner och rader  
När Du vill flytta rader och kolumner använder Du Alt-tangenten som startsignal.  
När Du använder Alt-tangenten i kombination med motsvarande piltangent förminskar / förstorar Du hela raden / kolumnen i tabellen med utgångspunkt från den högra / nedre kanten.  
Den högra / nedre kanten används som referenskant när Du håller ned skifttangenten.  
Om Du endast vill flytta den markerade raden / kolumnen, så håller Du Ctrl-tangenten nedtryckt.  
Hur tabellen respektive kolumnerna / raderna uppför sig när Du flyttar dem beror på vilket läge Du väljer.  
Om Du t ex vill förstora en kolumn utan att övriga kolumners kolumnbredd påverkas, väljer Du alternativet variabel.  
Infoga och radera kolumner och rader  
Om Du snabbt och enkelt vill infoga / ta bort en kolumn / rad i den aktuella tabellen, så aktiverar Du denna funktion genom att hålla ned Alt-tangenten tillsammans med Insert - eller Delete-tangenten.  
Det valda läget är nu aktiverat under cirka 3 sekunder (efter det att Du har släppt upp båda tangenterna).  
Inom denna tidsperiod kan Du trycka på den pilknapp i vars riktning den rad / kolumn befinner sig som ska infogas / tas bort.  
När Du har använt funktionen eller när tidsperioden har gått ut, upphävs det aktiverade läget.  
Hur tabeller uppför sig i textdokument, definierar Du i Verktyg - Alternativ... - Textdokument - Tabell.  
Textflöde  
Här kan du bland annat definiera textflödet i texten före och efter tabellen.  
Textflöde  
I det här området väljer du inställningar för textflödet före och efter tabellen.  
Du definierar typ av brytning, sidformatmallen som ska användas och upprepningen av tabellöverskriften.  
Brytning  
Med den här rutan aktiverar du tabellbrytningen.  
Välj typ av brytning från följande alternativfält:  
Sida  
Om du markerar det här alternativfältet infogas alltid en sidbrytning före eller efter tabellen.  
Om du bara vill undvika en sidbrytning inom tabellen, kan du markera hela tabellen och sedan klicka på ikonen Infoga - Ram på verktygslisten.  
Tabellen får en ram vars kant du kan ta bort via snabbmenyn på fliken Inramning.  
Nu kan tabellen inte längre brytas, men den kan heller inte bli längre än en sida.  
Kolumn  
Om Du markerar det här alternativfältet infogas alltid en kolumnbrytning före eller efter tabellen.  
Före  
Om Du markerar det här alternativet infogas sid - eller kolumnbrytningen före tabellen, och tabellen visas i början av nästa sida eller kolumn.  
Efter  
Om Du markerar det här alternativet infogas sid - eller kolumnbrytningen efter tabellen, och följande stycke visas i början av nästa sida eller kolumn.  
med sidformatmall  
Markera den här kryssrutan, om Du vill använda en viss sidmall efter sidbrytningen.  
Sidformatmall  
Välj önskad sidformatmall här.  
Sidnummer  
Om den automatiska sidnumreringen ska ändras på sidan efter sidbrytningen, anger Du önskat nummer för sidan som följer.  
Dela inte tabell  
Om Du vill förhindra en delning, måste Du markera den här kryssrutan.  
Håll ihop med följande stycke  
Om Du markerar den här kryssrutan hålls stycken ihop.  
Upprepa överskrift  
Markera den här rutan om du vill att innehållet på den första tabellraden ska användas som överskrift på den nya sidan efter en sidbrytning i tabellen.  
Om den här funktionen har valts, skrivs taggarna THEAD och TBODY vid export i HTML-format.  
Vertikal justering  
I det här området definierar Du den vertikala justeringen för texten i en cell.  
Överst  
Klicka på det här alternativet, om texten ska justeras vid cellens övre kant.  
Mitten  
Klicka på det här alternativet, om texten ska justeras i mitten av cellen.  
Underst  
Genom att klicka på det här alternativet justerar Du texten vid cellens nedre kant.  
Cell  
Det här kommandot är bara tillgängligt om du har markerat en tabell i dokumentet eller om markören står i en tabell.  
När Du har valt menykommandot Cell visas en undermeny med följande poster, som gäller enskilda celler i tabellen:  
Dela...  
Förbinda  
Här sammanfogas de markerade tabellcellerna till en cell.  
På det här sättet kan du exempelvis placera en huvudrubrik över två tabellkolumner.  
Det leder till felaktiga räkneresultat.  
Korrigera alla formler i tabellen när du har förbundit cellerna.  
Dela celler  
Här delar du en cell eller ett cellområde i ytterligare tabellceller.  
Dela  
Ange här antalet uppdelningar av den aktuella cellen eller det markerade cellområdet.  
Riktning  
Här anger Du om ytterligare kolumner eller rader ska infogas.  
horisontellt  
Ytterligare tabellrader infogas i den aktuella cellen eller det markerade cellområdet.  
vertikalt  
Ytterligare tabellkolumner infogas i den aktuella cellen eller det markerade cellområdet.  
Skydda  
Med det här kommandot skyddar du innehållet i markerade celler i en tabell.  
På så sätt ser du till att innehållet inte ändras eller raderas av misstag.  
Motsvarande kommandon är därför inte tillgängliga.  
Du kan däremot placera markören i ett skyddat cellområde och markera innehållet och t.ex. kopiera det.  
Om markören står i ett skrivskyddat cellområde visas detta med en upplysning på statuslisten.  
Om du vill upphäva cellskyddet, markerar du cellen resp. cellerna och väljer Format - Cell - Upphäv skydd.  
Upphäv skydd  
Med det här kommandot upphäver du cellskyddet för alla celler i den aktuella tabellen.  
Markören kan då stå i en skyddad cell eller i ett markerat område i tabellen.  
Det finns andra möjligheter att upphäva cellskyddet.  
Du kan upphäva skyddet för flera tabeller samtidigt genom att markera dem och sedan trycka på tangentkombinationen Kommando Ctrl +Skift+T.  
Även om markören står någonstans i dokumentet, dvs inte alls har någon förbindelse med någon cell eller tabell, kan Du upphäva cellskyddet för alla befintliga tabeller.  
Även här använder Du kortkommandot Kommando Ctrl +Skift+T.  
Du kan även nå funktionen för att upphäva cellskyddet från Navigator.  
Överst  
Det här kommandot är bara meningsfullt om cellen är större än vad texten i cellen kräver, om du t.ex. har anpassat cellens storlek fritt.  
Mitten  
Det här kommandot är bara meningsfullt om cellen är större än vad texten i cellen kräver, om du t.ex. har anpassat cellens storlek fritt.  
Underst  
Det här kommandot är bara meningsfullt om cellen är större än vad texten i cellen kräver, om du t.ex. har anpassat cellens storlek fritt.  
Rad  
Om du väljer det här menykommandot öppnas en undermeny med kommandon som gäller raderna i en tabell.  
Den här undermenyn är till för att ställa in radhöjd och för att markera, infoga och radera rader.  
Höjd  
Optimal höjd  
Infoga  
Radhöjd  
Med den här funktionen kan Du definiera en fast radhöjd.  
Denna höjd kan gälla för en tabellrad eller alla markerade tabellrader.  
Höjd  
Ange här önskad höjd för den aktuella tabellraden eller det markerade tabellområdet.  
anpassa dynamiskt  
Om Du markerar den här kryssrutan, anpassas radens höjd automatiskt till innehållets storlek.  
Om Du har ställt in höjden manuellt, anpassas inte tabellradens höjd till den text som Du matar in.  
Om Du vill återvända till den automatiska anpassningen, väljer Du Format - Rad - Optimal höjd.  
Optimal höjd  
Med det här kommandot anpassar du automatiskt tabellradens höjd till textinnehållet.  
Detta är standardinställningen för nya tabeller.  
Det här menyalternativet kan du bara använda om du har definierat en fast höjd för en tabellrad.  
Markera  
Med det här kommandot markerar du hela raden där markören står i tabellen.  
Det här menykommandot visas bara när markören står i en tabell.  
Radera  
Med hjälp av den här funktionen raderar du den aktuella tabellraden.  
Du ombeds inte bekräfta raderingen.  
De följande tabellraderna flyttas en position uppåt.  
Fördela raderna jämnt  
Med det här kommandot blir höjden för de markerade raderna identisk.  
Då tilldelas alla rader den största radhöjden.  
Kolumn  
Till det här menykommandot hör en undermeny med kommandon som gäller kolumnerna i den aktuella tabellen.  
Där finns kommandon för att ställa in kolumnbredd och markera, infoga och radera kolumner.  
Kommandot Kolumn visas bara när textmarkören står i en tabell.  
Bredd...  
Optimal bredd  
Infoga...  
Kolumnbredd  
Med den här funktionen ändrar du bredden på de markerade kolumnerna i tabellen.  
Det här menykommandot är bara tillgängligt när markören står i en tabell.  
Bredd  
Här ställer Du in kolumnbredden för en enskild kolumn.  
Kolumn  
Här anger Du numret på den kolumn som ska ändras, eller också använder Du mallen för den aktuella kolumnen.  
Bredd  
Ange här den önskade kolumnbredden.  
När Du ändrar en kolumnbredd gäller detta alltid även bredden på följande kolumn.  
När Du ändrar den sista kolumnen påverkas den första tabellkolumnen.  
Optimal bredd  
Med det här kommandot anpassas kolumnbredden till cellinnehållet.  
Ändringen av en kolumnbredd påverkar inte bredden på de andra tabellkolumnerna.  
Tabellen blir totalt inte bredare än vad sidbredden tillåter.  
Detta menykommando visas bara när markören står i en tabell.  
Markera  
Med det här kommandot markerar du hela kolumnen där markören står i tabellen.  
Det här menykommandot visas bara när markören står i en tabell.  
Infoga kolumner / rader  
Med den här funktionen kan du infoga kolumner resp. rader i en tabell.  
Det här menykommandot visas bara när markören står i en tabell.  
Infoga  
Här anger du det antal kolumner resp. rader som ska infogas.  
Position  
Här anger du placeringen av de kolumner resp. rader som ska infogas.  
framför  
Nya tabellrader infogas ovanför den aktuella raden eller det markerade området.  
bakom  
Ny tabellrader infogas under den aktuella raden eller det markerade området.  
Radera  
Med den här funktionen raderar du den aktuella tabellkolumnen.  
Du ombeds inte att bekräfta raderingen.  
De följande kolumnerna i tabellen flyttas ett steg åt vänster.  
Det här menykommandot visas bara när markören står i en tabell.  
Fördela kolumnerna jämnt  
Med det här kommandot tilldelas de markerade kolumnerna identisk bredd.  
Den totala bredden för alla kolumner adderas och fördelas på antalet markerade kolumner.  
Mallkatalog  
I mallkatalogen redigerar och organiserar du formatmallarna.  
Här kan du skapa, ändra, välja ut och organisera mallarna som används i det aktuella dokumentet.  
Alla inställningar i den här dialogrutan räknas som indirekt formatering.  
Förutom förvaltningen av mallar har Stylist samma funktionalitet.  
Om du vill göra ett dokument till en mall (dokumentmall), använder du kommandot Arkiv - Dokumentmall - Spara.  
Malltyp  
I mallkatalogen visas det aktuella områdets malltyp i en listruta.  
Om markören t.ex. står i ett textstycke visas styckeformatmallarna; om en ram är markerad visas ramformatmallarna.  
Klicka i listrutan om du vill välja en annan malltyp.  
Namn  
Betydelse  
Teckenformatmallar  
Teckenformatmallar används för indirekt formatering av enskilda tecken, ord eller meningar.  
Du kan även välja att t.ex. använda en viss teckenformatmall för ett ord i en text och en annan teckenformatmall för den omgivande texten.  
Styckeformatmallar  
Styckeformatmallar används för indirekt formatering av hela stycken.  
Förutom normala inställningar för styckeformatering innehåller styckeformatmallarna även information om vilket teckensnitt används i stycket och nästa formatmall.  
Ramformatmallar  
Ramformatmallar används för indirekt formatering av grafik - och textramar.  
Genom att använda ramformatmallar sparar du tid, eftersom grafikobjekten och ramarna då automatiskt får önskat format.  
Sidformatmallar  
Sidformatmallar används för indirekt formatering av hela sidor.  
När du definierar formatmall för följande sida ser %PRODUCTNAME till att den nya sidan får definierat sidformat vid automatisk sidbrytning.  
Numreringsformatmallar  
Numreringsformatmallar används för formatering av stycken i numreringar eller punktuppställningar.  
Mallista  
Den som för tillfället används är markerad.  
Om du vill redigera en mall använder du snabbmenyn och om du vill tilldela en mall dubbelklickar du på den.  
På snabbmenyn kan du välja kommandon för att skapa en ny mall, radera en mall som du själv har skapat eller ändra den markerade mallen.  
Mallområde  
För att förteckningen ska bli överskådlig är mallarna uppdelade i olika mallområden.  
Välj ett annat mallområde för den aktuella malltypen om den önskade mallen inte finns på listan.  
Namn  
Betydelse  
Automatiskt  
Visar de mallar som passar i det aktuella sammanhanget.  
Alla formatmallar  
Visar alla mallar av den aktuella malltypen.  
Använda formatmallar  
Visar de mallar av den aktuella malltypen som används i det aktuella dokumentet.  
Du kan även välja dem på objektlisten.  
Användardefinierade formatmallar  
Visar de användardefinierade mallarna av den aktuella malltypen.  
Textformatmallar  
Visar de mallar som kan användas för text.  
Kapitelformatmallar  
Visar de mallar som kan användas för kapitel.  
Listformatmallar  
Visar de punktuppställnings - och numreringsformatmallar som kan användas för listor.  
Förteckningsformatmallar  
Visar de mallar som kan användas för förteckningar.  
Formatmallar specialområde  
Visar mallar som kan användas i särskilda områden (t.ex. sidhuvuden, fotnoter, tabeller, bildtexter).  
HTML-formatmallar  
Visar mallar för HTML-dokument.  
Villkorliga mallar  
Visar de mallar för vilkas användning Du har definierat villkor.  
Hierarkiskt  
Visar mallarna i den aktuella malltypen i en hierarkisk uppställning.  
Den här visningen liknar visningen av hårddiskens mappstruktur.  
Om Du vill se mallarna på en underliggande nivå klickar Du på plustecknet intill mallnamnet.  
Nytt...  
Klicka på den här kommandoknappen om du vill skapa en ny mall.  
Alltefter vald malltyp visas dialogrutan Styckeformatmall, Teckenformatmall, Ramformatmall, Sidformatmall eller Numreringsformatmall.  
Ändra...  
Klicka på den här kommandoknappen om Du vill ändra den mall som är markerad i listrutan eller vill undersöka inställningarna i den aktuella mallen.  
Motsvarande malldialogruta öppnas.  
Radera...  
Du blir först ombedd att bekräfta.  
Du kan bara radera användardefinierade mallar.  
Administrera...  
Klicka på den här kommandoknappen när Du vill kopiera de mallar som används i det aktuella dokument till andra dokument, eller omvänt kopiera mallar från andra dokument till det aktuella dokumentet.  
Dialogrutan Administrera dokumentmallar öppnas.  
Styckeformatmall  
Här skapar eller ändrar du en styckeformatmall.  
Fliken Villkor visas bara om du skapar en ny styckeformatmall eller om du ändrar en villkorlig mall.  
Om du ändrar en mall, som inte är en villkorlig mall, visas inte den här fliken.  
Teckenformatmall  
Här kan du skapa en teckenformatmall.  
Ramformatmall  
Här kan du skapa en ramformatmall.  
Numreringsformatmall  
Här kan du skapa en numreringsformatmall.  
Numreringsformatmallar förvaltas i Mallkatalogen och är tillgängliga i Stylist där du kan använda dem för att utforma dokumentet.  
När en numreringsformatmall skapas tilldelas numreringen ett namn, därför kallas sådana formatmallar namngivna numreringar.  
Ej namngivna numreringar, som används för direkt formatering, kan du skapa med dialogrutan Numrering / punktuppställning eller med ikonerna på objektlisten för punktuppställningar och numreringar.  
Villkor  
Här kan du definiera villkoren för villkorliga formatmallar.  
När du definierar en ny mall kan du ange om den ska vara "villkorlig".  
Däremot kan du ändra själva villkoren.  
Om det stycke som har formaterats med en villkorlig mall står i ett sammanhang som är kopplat till en använd mall, används den styckeformatmall som hör till sammanhanget.  
Om ingen mall har kopplats till sammanhanget, gäller de attribut som är definierade i den villkorliga mallen.  
Följande exempel förtydligar det här sambandet:  
Öppna ett tomt textdokument och skriv ett kort affärsbrev med ett brevhuvud (Format - Sida... - Sidhuvud).  
Definiera en ny styckeformatmall genom att ge kommandot Nytt... på snabbmenyn till Stylist för styckeformatmallar och ange alla styckeegenskaper som Du vill att normala stycken i affärsbrevet ska ha i dialogrutan Styckeformatmall.  
Döp mallen till "Affärsbrev".  
På det sättet definierar Du den nya styckeformatmallen som villkorlig mall.  
Välj posten Sidhuvud under Sammanhang, och välj den mall som ska gälla för sidhuvudena i affärsbrevet, t ex den fördefinierade styckeformatmallen "Sidhuvud" i listrutan Styckeformatmallar. (Naturligtvis kan Du här välja en mall som Du själv har definierat.)  
Genom att dubbelklicka på den valda posten i listrutan Styckeformatmallar, eller genom att klicka på Tilldela, tilldelar Du styckeformatmallen det nya sammanhanget.  
Stäng nu dialogrutan för styckeformatmallar med OK och formatera alla stycken i affärsbrevet inklusive sidhuvudet med den nya, villkorliga styckeformatmallen "Affärsbrev". (När Du klickar i sidhuvudet kan Du i förekommande fall behöva ta fram alla mallar eller användarmallar i Stylist för att kunna använda den nya mallen "Affärsbrev".)  
Du ser nu att texten i sidhuvudet har de attribut som har definierats i styckeformatmallen "Sidhuvud" (om det var den Du använde), medan alla andra delar av dokumentet har de attribut som Du definierade i den (villkorliga) styckeformatmallen "Affärsbrev ".  
Vi har skapat mallen "Brödtext" som villkorlig mall.  
Alla mallar som du själv skapar och baserar på "Brödtext" kan därför också användas som villkorliga mallar.  
När Du exporterar till ett annat format (RTF, HTML osv) skrivs den styckeformatmall som har tilldelats sammanhanget.  
som villkorlig mall  
Markera detta fält när Du definierar en ny mall, om Du vill att den nya mallen ska vara en villkorlig mall.  
Sammanhang  
Disposition nivå 1 - 10, Numrering / punktuppställning nivå 1 - 10, Tabellhuvudrad, Tabellinnehåll, Område, Ram, Fotnot, Sidhuvud och Sidfot.  
Använda formatmallar  
Här visas en lista över alla styckeformatmallar som har tilldelats ett visst sammanhang.  
Styckeformatmallar  
I listrutan visas en lista över alla styckeformatmallar som Du kan tilldela ett visst sammanhang.  
Ta bort  
Klicka här om Du vill ta bort den markerade tilldelningen av sammanhang och använd mall.  
Tilldela  
Om Du klickar på kommandoknappen Tilldela, tilldelas den markerade styckeformatmallen det tidigare valda sammanhanget som använd mall.  
Stylist  
Med Stylist tilldelar du objekt och textområden mallar.  
Du uppdaterar mallarna, ändrar befintliga mallar och skapar nya mallar.  
Stylists förankringsbara fönster kan vara öppet medan du redigerar dokumentet.  
Uppe i Stylist-fönstret finns ikoner för formatering av dokument:  
Malltyper  
Styckeformatmallar  
Den här ikonen visar Styckeformatmallarna i Stylist-fönstret.  
Styckeformatmallar används för mjuk formatering av hela stycken.  
Teckenformatmallar  
Den här ikonen visar Teckenformatmallarna i Stylist-fönstret.  
Teckenformatmallar används för indirekt formatering av enskilda tecken, ord eller meningar.  
Ramformatmallar  
Den här ikonen visar Ramformatmallarna i Stylist-fönstret.  
Ramformatmallar används för mjuk formatering av grafik - och textramar.  
Sidformatmallar  
Den här ikonen visar Sidformatmallarna i Stylist-fönstret.  
Sidformatmallar används för mjuk formatering av sidstrukturen.  
Numreringsformatmallar  
Den här ikonen visar Numreringsformatmallarna i Stylist-fönstret.  
Numreringsformatmallar används för indirekt formatering av numreringar och punktuppställningar.  
Tilldelningsläge  
Med den här ikonen växlar du till ett läge där du kan använda den aktuella formatmallen på objekt och texter med musen.  
När du vill lämna tilldelningsläget klickar du en gång till på ikonen eller trycker på Esc.  
Ny formatmall av markering  
Den får det markerade styckets, objektets eller tecknets format.  
Du ger den nya mallen ett namn i dialogrutan Skapa formatmall.  
Uppdatera formatmall  
Om du klickar på den här ikonen ersätts styckeformatmallen som är markerad i Stylist med formateringen som det markerade stycket har.  
Mallista / Mallområde / Snabbmeny Nytt... / Ändra... / Radera...  
I Stylist har du tillgång till samma funktioner som i dialogrutan Mallkatalog.  
Använda formatmallar  
AutoFormat  
Här kan du bearbeta textdokument automatiskt enligt vissa regler.  
Reglerna definierar du under Verktyg - AutoKorrigering.  
När textmarkören står i en tabell visas dialogrutan AutoFormat om du väljer kommandot AutoFormat.  
Under inmatningen  
Alternativen för AutoFormat ställer du in under fliken Alternativ i dialogrutan AutoKorrigering, som du öppnar med kommandot Verktyg - AutoKorrigering / AutoFormat...  
Du kan använda AutoFormat för formatering av textdokument och ren ASCII-text.  
Du kan inte ändra hårda teckenformateringar med AutoFormat.  
Ordkompletteringar sker redan medan Du skriver, förutsatt att Du redan har skrivit ordet en gång, så att den automatiska korrigeringen kan hämta det ur "minnet".  
Ytterligare regler för AutoFormat  
Om den automatiska formateringen inte passar, kan Du ångra den direkt med kommandot Ångra.  
AutoFormat för tabeller  
Med AutoFormat formateras tabellen automatiskt.  
Så formaterar du en tabell automatiskt  
Placera markören i en valfri cell i texttabellen eller markera några celler.  
Välj kommandot AutoFormat på menyn Format och välj ett format.  
Klicka på OK.  
Cellformat  
I den här listrutan visas ett urval av fördefinierade format.  
Lägg till  
Här lägger du till ett nytt AutoFormat på listan.  
Gör så här:  
Formatera en tabell i önskat format.  
Markera den och öppna dialogrutan AutoFormat.  
Klicka på kommandoknappen Lägg till.  
Ange ett namn på det nya AutoFormatet i nästa dialogruta, Lägg till AutoFormat.  
Radera  
Med den här kommandoknappen raderar du, efter att ha bekräftat detta i en dialogruta, det markerade AutoFormatet från listan.  
Fler  
Med den här kommandoknappen utvidgar du.  
Du stänger tilläggsområdet i dialogrutan genom att klicka en gång till.  
Formatering  
Avmarkera här den formatering som inte ska skapas automatiskt.  
Talformat  
Markera här om om talformatet ska inkluderas i AutoFormatet.  
Teckensnitt  
Markera här om teckensnittet ska inkluderas i AutoFormatet.  
Justering  
Markera här om cellinnehållets justering ska användas.  
Inramning  
Markera här om stilen för inramning av celler ska användas.  
Mönster  
Markera här om bakgrundsmönstret ska inkluderas i AutoFormatet.  
Byt namn  
Här döper du om en markerad post i listan Cellformat.  
Kombinera  
Minsta storlek  
I detta rotationsfält definierar Du hur breda (i procent av den skrivbara sidbredden) enradiga stycken minst måste vara för att de automatiskt ska kombineras till ett enda stycke.  
Använd  
Med det här kommandot startar du den automatiska formateringen (i efterhand) av hela det aktuella textdokumentet.  
För automatisk formatering gäller följande regler:  
AutoFormat för överskrifter  
Ett stycke formateras som överskrift om det finns ett tomt stycke ovanför och nedanför, om raden börjar med en stor bokstav och om den inte avslutas med punkt (.), komma (,) eller semikolon (;).  
Överskriftsnivåerna bestäms av antalet blanksteg eller tabbtecken.  
Om Du placerar ett blanksteg i början av raden, formateras överskriften på den högsta nivån.  
Om Du placerar ett tabbtecken i början av raden, blir det likaså en överskrift på den högsta nivån; två tabbtecken ger en överskrift på nivå två osv.  
Ett kolon sist på raden ger likaså en överskrift på nivå tre.  
När respektive format har tilldelats överskriften, tas det följande tomma stycket bort, och nästa stycke får det format som är inställt som Nästa formatmall.  
AutoFormat för numrering / punktuppställning  
Om du inleder ett stycke med ett bindestreck (-), en asterisk (*) eller ett plustecken (+), eller med ett tvåställigt tal och ett blanksteg eller ett tabbtecken, formateras en punktuppställning / numrering som du därefter kan redigera.  
När det gäller tal inkluderas de tecken som står före eller efter punktuppställningen / numreringen i formateringsregeln.  
Respektive nivå bestäms av talet / avgränsaren.  
Den automatiska numreringen aktiveras bara i stycken som formaterats med någon av styckeformatmallarna "Standard", "Brödtext" eller "Brödtext indrag ".  
Autoformat för skiljelinjer  
Om Du gör ett stycke som består av minst tre bindestreck (-- -), understreck (___) eller likhetstecken (===), ersätts det av en skiljelinje med en längd lika med sidans bredd.  
Linjen skapas som undre inramning av föregående stycke.  
Därvid gäller följande:  
Bindestreck (-) ger en enkel linje, 0,05 punkter tjock och med avståndet 0,75 mm.  
Understreck (_) ger en enkel linje, 1 punkt tjock och med avståndet 0,75 mm.  
Likhetstecken (=) ger en dubbel linje, 1,10 punkter tjock och med avståndet 0,75 mm.  
Använd och redigera ändringar  
Med det här kommandot startar du den automatiska formateringen i hela det aktuella textdokumentet.  
Du kan redigera ändringarna i efterhand.  
Kommandot öppnar en dialogruta med tre kommandoknappar, med vars hjälp Du i efterhand kan bestämma vad som ska hända med ändringarna.  
Acceptera alla  
Med Acceptera alla accepterar Du alla ändringar Du gjort.  
Avböj allt  
Om du klickar på den här kommandoknappen kastar du bort alla ändringar.  
Redigera ändringar  
Med den här kommandoknappen öppnar du dialogrutan Acceptera eller ignorera Autoformat-ändringar.  
Under fliken Lista kan du ignorera resp. acceptera enstaka ändringar.  
Om du vill se ändringar som en viss författare har gjort eller ändringarna under en viss tidsperiod, kan du ställa in det under fliken Filter.  
Ladda mallar  
Här laddar du formatmallar från ett annat dokument eller från en dokumentmall i det aktuella dokumentet.  
Kategorier  
Dokumentmallarna är indelade i kategorier efter innehåll.  
Här väljer du en kategori.  
Mallar  
Här väljer du en dokumentmall i den valda kategorin.  
Text  
Markera den här rutan om du vill använda textformatmallarna från det markerade dokumentet i det aktuella dokumentet.  
Till textmallarna hör stycke - och teckenformatmallarna.  
Ram  
Markera den här rutan om du vill använda ramformatmallarna från det markerade dokumentet i det aktuella dokumentet.  
Sidor  
Markera den här rutan om du vill använda sidformatmallarna från det markerade dokumentet i det aktuella dokumentet.  
Numrering  
Markera den här rutan om du vill använda numreringsformatmallarna från det markerade dokumentet i det aktuella dokumentet.  
Skriv över  
Markera den här rutan om formatmallarna i det aktuella dokumentet ska ersättas med det andra dokumentets mallar med samma namn.  
När befintliga formatmallar skrivs över sker det utan säkerhetskontroll.  
Från fil  
Här öppnar du en dialogruta för filurval där du kan ladda formatmallar från ett annat dokument.  
Textanpassning  
På undermenyn till Format - Textanpassning bestämmer du hur en text ska förhålla sig till ramar, grafikobjekt och objekt.  
Ingen textanpassning  
Textanpassning sida  
Dynamisk textanpassning sida  
Textgenomflöde  
I bakgrunden  
Kontur  
Redigera kontur...  
Första stycket  
Redigera...  
Dela upp tabell  
Det här kommandot delar upp den aktuella tabellen i två tabeller vid cellmarkörens position.  
I en dialogruta kan du välja alternativ för uppdelningen.  
Samma kommando finns på snabbmenyn till tabeller i %PRODUCTNAME Writer.  
Läge  
Här väljer Du tabelluppdelningsläge.  
Kopiera överskrift  
Den första raden i utgångstabellen kopieras som extra första rad i den andra tabellen.  
Egen överskrift, med formatmall  
Den andra tabellen får en ny tom rad med formatmallen från den första raden i utgångstabellen.  
Egen överskrift  
Den andra tabellen får en ny tom rad.  
Ingen överskrift  
Tabellen delas utan ändringar.  
De kan bli ogiltiga vid delningen, vilket innebär att Du måste återskapa dem i efterhand.  
Förbinda tabell  
Med det här kommandot sammanfogar du två tabeller som står direkt efter varandra.  
Du kan också ångra delningen av en tabell med det här kommandot.  
Det här kommandot är bara tillgängligt, om de tabeller som ska sammanfogas står direkt efter varandra utan någon mellanliggande rad.  
Du raderar en tom rad med Delete-tangenten.  
Tabellraderna anpassas till varandra liksom de tabellformler som eventuellt ingår.  
Om tre tabeller står efter varandra och markören står i den mellersta när du förbinder tabellerna, öppnas en dialogruta där du tillfrågas med vilken av de båda den ska förbindas.  
Mallar  
Här har du tillgång till samtliga kommandon för hantering av mallar.  
Katalog...  
Ladda...  
Avstavning  
Med det här menykommandot aktiverar du avstavningen i %PRODUCTNAME Writer. %PRODUCTNAME Writer söker igenom dokumentet med avseende på om avstavning ska göras i radsluten.  
Om ett ord för eventuell avstavning påträffas, visar %PRODUCTNAME Writer en dialogruta där du kan bekräfta avstavningsstället eller korrigera det.  
Standardinställningarna för automatisk avstavning i %PRODUCTNAME Writer kan du ställa in under fliken Textflöde.  
Fliken finns i dialogen Stycke som Du öppnar genom att välja Format - Stycke.  
Om du vill redigera styckeformatmallen öppnar du snabbmenyn till ett stycke som har den här mallen och väljer där kommandot Redigera styckeformatmall.  
Träffarna visas i en dialogruta.  
Om du vill:  
Gör du så här:  
Bekräfta alla markerade avstavningar  
Klicka på Avstava  
Bekräfta en avstavningsposition som är utmärkt med =.  
Välj avstavning genom att markera den, eller genom att hoppa mellan avstavningsförslagen med hjälp av pilknapparna, och klicka på Avstava.  
Inte avstava ordet  
Klicka på Ta bort  
Avbryta hela funktionen  
Klicka på Avbryt  
Med Kommando Ctrl +minustecken skriver du ett användardefinierat bindestreck.  
Om du tycker att visningen av bindestreck mitt i raderna stör, väljer du Verktyg - Alternativ - Textdokument - Formateringshjälp och avmarkerar rutan Användardefinierade bindestreck.  
Ett skyddat bindestreck förbinder två orddelar som inte får delas sist på en rad.  
För att du ska kunna göra det måste du öppna dialogen Anpassa via Verktyg - Anpassa... och koppla funktionen "Infoga hårt bindestreck" till en tangent i funktionsområdet "Infoga ".  
Det finns ett exempel på hur en funktion kopplas till en tangent i > %PRODUCTNAME -hjälpen.  
Avstavningen genomförs utan att du tillfrågas om du aktiverar alternativet Automatisk avstavning under Verktyg - Alternativ - Språkinställningar - Lingvistik.  
Om du vill utesluta enskilda stycken från den automatiska avstavningen, markerar du dem som block, väljer kommandot Format - Stycke och klickar på fliken Textflöde där du avmarkerar alternativet Automatisk i området Avstavning.  
Ord  
I det här området hittar du textfältet Ord.  
Ord  
Här visas det ord som ska avstavas.  
Du kan ta bort dem och infoga nya.  
Höger / vänsterpil  
Om det finns flera avstavningsmöjligheter i ordet, kan du flytta mellan dem med pilknapparna.  
Nästa  
Klicka här om ordet inte ska avstavas men avstavningskontrollen ska fortsätta.  
Avstava  
Klicka här om ordet ska avstavas på angiven plats.  
Ta bort  
Klicka här om du inte vill avstava ett ord.  
Alla visade avstavningsställen i ordet tas bort i den här avstavningsgenomgången; även de som du har ställt in manuellt med Kommando Ctrl och bindestreck.  
Kapitelnumrering  
Med den här funktionen definierar du kapitelnumreringens typ och utseende.  
De här inställningarna gäller för det aktuella dokumentet.  
En kapitelnumrering är kopplad till en styckeformatmall.  
Om du definierar en kapitelnumrering för en styckeformatmall, t.ex. "Överskrift1", används den numreringen alltid när mallen används.  
Du kan definiera upp till 10 kapitelnivåer och skapa olika numreringar för olika nivåer.  
Definitionen för varje enskild nivå anger du i dialogrutan Kapitelnumrering.  
Kapitelnumreringarna visas med grå bakgrund i dokumentet om du aktiverar kommandot Markeringar på menyn Visa.  
Format  
Om du klickar på den här kommandoknappen, kan du spara den inställda kapitelnumreringsdefinitionen eller välja en redan definierad och sparad kapitelnumrering på popupmenyn.  
Medan en kapitelnumrering, som du har definierat i dialogrutan Kapitelnumrering, är kopplad till det aktuella dokumentet, har du tillgång till sparade definitioner för kapitelnumreringar i alla textdokument.  
Kommandoknappen Format visas bara för kapitelnumrering.  
För numreringar eller punktuppställningar av enskilda stycken kan du arbeta med numreringsformatmallar, så att du alltid har tillgång till numreringen eller punktuppställningen om du definierar den som mall.  
Namnlös 1 - 9  
Genom att välja någon av de här posterna tilldelar Du den aktuella numreringsnivån ett fördefinierat numreringsformat.  
På popup-menyn visas som standard nio olika poster, till en början med de förinställda namnen "Namnlös 1" t o m "Namnlös 9 ".  
Du kan ersätta dem med egna inställningar och namn i den dialogruta som Du öppnar med kommandot Spara som....  
Spara som...  
Med det här menykommandot öppnar Du en dialogruta för att spara ett kapitelnumreringsformat.  
Den kapitelnumrering som Du sparar på detta vis, kan Du när som helst använda genom att klicka på kommandoknappen Format på popup-menyn.  
Spara som  
Välj här den post i den undre listrutan som Du vill använda som namn på den kapitelnumrering som ska sparas.  
I den övre listrutan kan Du redigera den valda posten och ge kapitelnumreringen ett nytt namn.  
Klicka sedan på OK.  
Namnet på kapitelnumreringen visas nu på popup-menyn, och på så vis har Du alltid tillgång till det.  
Numrering  
Här definierar du visningstyp för kapitelnumreringen.  
Nivå  
Här väljer du en kapitelnivå som du vill definiera en numrering för.  
Om du markerar en speciell nivå, visas de aktuella formateringsinställningarna och den använda styckeformatmallen i respektive fält på sidan under fliken.  
Med alternativet "1 - 10" kan du göra inställningar som ska gälla för alla kapitelnivåer.  
De är sedan inte knutna till en viss styckeformatmall.  
Numrering  
Här definierar du styckeformatmallen för kapitelnumreringen och bestämmer numreringstyp och skiljetecken.  
Styckeformatmall  
Klicka i fältet och välj önskad styckeformatmall för den markerade nivån.  
Det innebär att respektive kapitelnivå inte definieras.  
Nummer  
I det här kombinationsfältet väljer du numreringstyp för den eller de aktuella nivåerna.  
Urval  
Funktion  
A, B, C,...  
Versaler  
a, b, c,...  
Gemener  
I, II, III,...  
Versala romerska siffror  
i, ii, iii,...  
Gemena romerska siffror  
1, 2, 3,...  
Arabiska siffror  
A,...  
AA,...  
AAA,...  
Antalet bokstäver återspeglar kapitelnivån.  
Andra numreringen på tredje nivån blir alltså "BBB".  
a,... aa,... aaa,...  
Antalet bokstäver återspeglar kapitelnivån.  
Tredje numreringen på andra nivån blir alltså "cc".  
Utan  
Inga numreringstecken.  
Endast de tecken som har definierats som skiljetecken visas vid radens början.  
Teckenformatmall  
Markera här teckenformatmallen för numreringstecknet.  
Fullständig  
I det här rotationsfältet kan du ställa in hur många överordnade nivåer som ska visas för den eller de aktuella kapitelnivåerna.  
Du kan t.ex. visa numreringar på den tredje nivån i kapitel 2 som 2.1.1, 2.1.2, 2.1.3 och så vidare.  
Skiljetecken framför  
Om vissa tecken ska placeras framför numreringen anger du dem här.  
Med "Kapitel" får du exempelvis numreringen "Kapitel 1 ", om du använder arabiska siffror för numreringen.  
Skiljetecken bakom  
Om du vill infoga ytterligare ett eller flera tecken efter de automatiskt skapade numreringstecknen, så kan du ange dem här.  
Med "kapitlet" får du t.ex. numreringen "1 kapitlet ", om du använder arabiska siffror för numreringen.  
Börja med  
Här definierar du vilket nummer eller tecken som kapitelnumreringen ska börja med.  
Om du t.ex. har skapat ett nytt dokument för det andra kapitlet i ditt arbete, anger du här värdet 2 för den första kapitelnivån.  
Om du infogar en numrering eller punktuppställning inom ett stycke på en sida, d.v.s. i direkt anslutning till en text, tilldelas numreringen eller punktuppställningen stycket.  
Fotnotsinställning  
Här definierar du vilka fotnotsinställningar som ska användas.  
Det finns olika inställningsmöjligheter för fot - och slutnoter.  
De inställningar som du gör här är giltiga för hela textdokumentet.  
Fotnoter  
Den här fliken använder du för att utforma fotnoter.  
Du har tillgång till följande möjligheter: placering av fotnoterna i dokumentet, typ av fotnotsnumrering, val av formatmallar som ska användas och inmatning av hänvisningstexter.  
Funktioner för formatering av fotnotsområdet finns under menykommandot som beskrivs här, Verktyg - Fotnoter och under Format - Sida... - Fotnot.  
Automatisk numrering  
Här definierar du typ av fotnotsnumrering och vilken omfattning den ska ha.  
Numrering  
Här väljer du typ av numrering  
Urval  
Funktion  
A, B, C  
Stora bokstäver  
a, b, c  
Små bokstäver  
I, II, III  
Stora romerska siffror  
i, ii, iii  
Små romerska siffror  
1, 2, 3  
Arabiska siffror  
A,...  
AA,...  
AAA,...  
Alfabetisk numrering med likadana stora bokstäver.  
Men alla ytterligare numreringar förses därefter alltid med likadana bokstäver:  
Efter Z (26) följer AA (30), BB (31), CC (32) osv.  
a,... aa,... aaa,...  
Alfabetisk numrering med likadana små bokstäver.  
Efter z (26) följer aa (27), bb (28), cc (29) osv.  
Räkning  
Här definierar du om den automatiska fotnotsnumreringen ska göras fortlöpande per sida, per kapitel eller i hela dokumentet.  
När du ska ange numreringens giltighet har du följande alternativ:  
Alternativ  
Betydelse  
Per sida  
Alla fotnoter på en sida numreras fortlöpande, och på nästa sida börjar numreringen om igen. (Det här alternativet är bara tillgängligt om du har valt alternativet Sidslut under Placering.)  
Per kapitel  
Alla fotnoter i ett kapitel numreras fortlöpande, och i nästa kapitel börjar numreringen om.  
Per dokument  
Alla fotnoter i dokumentet numreras löpande.  
Börja med  
Om du väljer alternativet Per dokument för numreringen, kan du definiera med vilket fotnotsnummer numreringen ska börja här.  
Detta kan vara praktiskt om fotnotsnumreringen ska omfatta flera dokument.  
Framför  
Om du vill infoga ett eller flera tecken framför fotnotssymbolen anger du dem här.  
Med "Not" får du exempelvis fotnotspresentationen "Not 1 ", om du använder en numrering med arabiska siffror.  
Bakom  
Om du vill infoga ett eller flera tecken efter fotnotssymbolen anger du dem här.  
Med ")" får du exempelvis fotnotspresentationen "1) ", om du använder en numrering med arabiska siffror.  
Lägg märke till att dessa tecken, som infogas före eller efter fotnotssymbolen, bara används vid den automatiska numreringen.  
Placering  
Det val du gör här anger om fotnoterna ska placeras längst ned på varje sida eller samlas i slutet av dokumentet.  
Sidslut  
De fotnoter som hör till en sida placeras alltid längst ned på sidan.  
Dokumentslut  
Alla fotnoter i dokumentet samlas i dokumentets slut. (På så sätt blir fotnoterna i praktiken slutnoter.)  
Formatmallar  
Det är bäst att formatera fotnotstexten med hjälp av mallar så att alla fotnoter i dokumentet (eller dokumenten) får ett enhetligt utseende.  
På så vis kan du lätt göra ändringar i formateringen av alla fotnoter genom att ändra mallen.  
Stycke  
Här väljer du styckeformatmallen för fotnotstexten.  
Det finns en fördefinierad styckeformatmall för fotnoter i förinställningen. %PRODUCTNAME har dessutom fler styckeformatmallar.  
När du ska ställa in en egen styckeformatmall för fotnoter här, öppnar du Stylist och definierar mallen under "Formatmallar specialområden".  
De förs sedan in i kombinationsfältet under fliken Fotnoter.  
Sida  
Här väljer du sidformatmall för fotnoter som ska samlas i dokumentets slut.  
Det finns en fördefinierad sidformatmall för fotnoter som standard.  
Dessutom hittar du samtliga fördefinierade sidformatmallar här, såväl de formatmallar som %PRODUCTNAME tillhandahåller som de som du har definierat själv.  
Du kan bara välja en sidformatmall om du har markerat alternativfältet Dokumentslut under Placering.  
Teckenformatmallar  
I det här området kan du tilldela fotnotssymbolerna formatmallar.  
Alla definierade teckenformatmallar är tillgängliga, inklusive mallarna för fotnotsankare och -tecken.  
Du kan använda de föreslagna teckenformatmallarna eller formatera fotnotssymbolerna med andra mallar som du vill.  
Textområde  
Välj önskad formatmall för symbolen i dokumentets textområde från listan.  
Fotnotsområde  
Här väljer du teckenformatmall för symbolen för dokumentets fotnotsområde.  
Hänvisningstext för flersidiga fotnoter  
Här kan du definiera meddelandetexter som ska infogas som förtydliganden vid flersidiga fotnoter.  
Vid slutet av fotnoten  
Här anger du den text som talar om att fotnoten fortsätter på nästa sida, t.ex. "Forts. på nästa sida". %PRODUCTNAME Writer lägger automatiskt till sidnumren till texten.  
På följande sida  
Här anger du den text som talar om att det rör sig om en fortsättning av fotnoterna från föregåande sida, t.ex. "Forts. från sida". %PRODUCTNAME Writer lägger automatiskt till sidnumren till texten.  
Slutnoter  
Här kan du utforma slutnoter.  
Du har tillgång till följande möjligheter: typ av slutnotsnumrering och val av de mallar som ska användas.  
Automatisk numrering  
Börja med  
Här kan du definiera med vilket slutnotsnummer numreringen ska börja.  
Det här är en användbar funktion om slutnotsnumreringen ska löpa genom flera dokument.  
Framför  
Om du vill infoga ett eller flera tecken framför slutnotssymbolen, så kan du skriva in dem här.  
Med "till" får du t.ex. slutnotsvisningen "till 1 "om du använder numrering med arabiska siffror.  
Bakom  
Om du vill infoga ett eller flera tecken efter slutnotssymbolen, så kan du skriva in dem här.  
Med ")" får du t.ex. slutnotsvisningen "1) "om du använder numrering med arabiska siffror.  
Observera att dessa tecken som ska infogas som tillägg framför eller bakom slutnotssymbolen bara används vid automatisk numrering.  
Formatmallar  
Du bör helst formatera slutnotstexten med hjälp av formatmallar, så att alla slutnoter i dokumentet (eller dokumenten) får ett enhetligt utseende.  
På så vis kan du lätt ändra formateringen för alla slutnoter genom att ändra formatmallen.  
Stycke  
Här väljer du styckeformatmall för slutnotstexten.  
Om du vill kunna ställa in en egen styckeformatmall för slutnoter här, öppnar du Stylist och definierar formatmallen under "Formatmallar specialområde".  
Mallen finns sedan med i kombinationsfältet under fliken Slutnoter.  
Sida  
Här väljer du sidformatmall för slutnoter.  
Förinställningen innehåller en fördefinierad sidformatmall för slutnoter.  
Dessutom hittar du samtliga fördefinierade sidformatmallar här, såväl de formatmallar som %PRODUCTNAME tillhandahåller som de som du har definierat själv.  
Teckenformatmallar  
I det här området kan du tilldela dokumentets slutnotssymboler formatmallar.  
Du kan välja bland alla definierade teckenformatmallar.  
Bland dessa finns formatmallarna slutnotsankare och -tecken.  
Du kan använda de föreslagna formatmallarna eller formatera slutnotssymbolerna som du vill med hjälp av andra formatmallar.  
Textområde  
Välj önskad formatmall för symbolen i dokumentets textområde i listan.  
Slutnotsområde  
Här väljer du teckenformatmall för slutnotssymbolen.  
Omvandla text till tabell  
Med den här funktionen omvandlar du en text till en tabell eller omvänt.  
Markera texten som ska göras om till en tabell, eller markera tabellen som ska göras om till text, och välj sedan det här kommandot.  
Dialogrutans utseende beror på i vilken riktning omvandlingen sker.  
Skiljetecken i text  
Här anger du vilket tecken som ska användas som skiljetecken.  
Varje styckeväxling i en text som ska omvandlas ger en ny rad i tabellen, och varje tabellrad utgör efter omvandling till text ett eget stycke.  
När du omvandlar en markerad tabell till normal text avgränsas innehållet i tabellens kolumner med det tecken som du väljer.  
Tabulator  
Tabbtecken gäller som skiljetecken.  
När du omvandlar text till tabell görs tabbpositionerna om till motsvarande kolumnbredder om du vill.  
Semikolon  
Semikolon (;) gäller som skiljetecken.  
Stycke  
%PRODUCTNAME skapar en tabell med en kolumn av texten.  
Varje stycke görs om till en tabellrad.  
Varje rad i tabellen blir ett eget stycke.  
Andra:  
Markera det här fältet när du vill ange ett annat skiljetecken än de alternativ som har beskrivits ovan.  
Som skiljetecken gäller det tecken som finns i textfältet intill.  
Textfält  
I det här fältet anger du vilket tecken som ska användas om du tidigare har aktiverat alternativfältet Andra.  
Samma bredd på alla kolumner  
Om du markerar det här fältet får alla kolumner i den nya tabellen samma kolumnbredd, oavsett var tabbtecknen står i texten.  
AutoFormat...  
Alternativ  
Här väljer du fler alternativ för omvandling från text till tabell.  
Överskrift  
Om du markerar den här rutan, formateras den första raden i den nya tabellen som överskrift.  
Upprepa på varje sida  
Om du markerar den här rutan, upprepas första raden i den nya tabellen på varje sida, om tabellen sträcker sig över flera sidor.  
Dela inte tabell  
Om du markerar den här rutan, placeras tabellen på en enda sida om det är möjligt.  
Inramning  
Om du markerar den här rutan, förses alla celler i den nya tabellen samt hela tabellen med en ram.  
Sortera  
Med det här kommandot sorterar du en markerad text radvis.  
Du kan definiera upp till tre sorteringsnycklar för sorteringen.  
Du kan kombinera alfanumeriska och numeriska sorteringsnycklar.  
Regel  
Nyckel 1 - 3  
Du använder de markerade nycklarna för sortering av de markerade områdena eller av tabellen.  
Du kan använda sorteringsnycklarna för sig eller i kombination.  
Kolumn 1 - 3  
Här anger du i vilken kolumn det ord står som ska användas som sorteringsvillkor.  
Tillåtet område är mellan 1 och 99.  
Om stycken ska sorteras bör du definiera vad som ska användas som avgränsningstecken under Avgränsare.  
Nyckeltyp 1 - 3  
Här anger du nyckeltyp.  
1, 12, 2.  
Ordning  
Raderna eller kolumnerna sorteras enligt 1, 2, 3 osv eller a, b, c osv.  
Fallande  
Raderna eller kolumnerna sorteras enligt 9, 8, 7 osv eller ö, ä, å osv.  
Riktning  
Kolumner  
Kolumnerna i en tabell sorteras efter den aktuella nyckeln.  
Rader  
Raderna i det markerade området eller tabellen sorteras efter den aktuella nyckeln.  
Avgränsare  
Stycken kan bara sorteras styckevis.  
Här kan du definiera avgränsare mellan stycken i listor.  
Tabulator  
Om de markerade styckena motsvarar en lista där styckena är avgränsade med tabbtecken, väljer du det här alternativet.  
Tecken  
Med hjälp av avgränsningstecknet kan %PRODUCTNAME bestämma positionen för sorteringsnycklarna (kolumnerna) i markerade stycken.  
...  
Den här kommandoknappen öppnar dialogrutan Specialtecken.  
Språk  
Välj språket, efter vars regler sorteringen sker, i det här fältet.  
Exakt jämförelse  
Om du aktiverar den här rutan genomförs en exakt jämförelse av stor och liten bokstav.  
Beräkna  
Med det här kommandot startar du beräkningen av formeln som finns i den aktuella markeringen.  
Resultatet lagras i urklippet.  
Sidformatering  
Med det här kommandot aktiverar du sidbrytningen av dokumentet manuellt. %PRODUCTNAME bryter automatiskt sidorna i dokumentet i bakgrunden.  
Aktuell status visas på statuslisten.  
När sidformateringen är klar, vilket kan ta en stund för mycket långa dokument, visas åter på statuslisten hur många sidor dokumentet omfattar totalt och på vilken sida markören står.  
Med det här kommandot ser du till att det sidantal som visas på statuslisten motsvarar dokumentets verkliga status.  
I normalfallet (vid "normallånga "dokument) bör detta automatiskt alltid vara fallet.  
När du arbetar med mycket långa dokument visas bara en uppskattning av sidantalet tills du väljer det här kommandot.  
Aktuell förteckning  
Med hjälp av det här kommandot kan du uppdatera den aktuella förteckningen.  
Förteckningen där markören står för tillfället, betraktas som aktuell förteckning.  
Om markören står i en förteckning hittar du förutom "Uppdatera förteckning" följande kommandon på snabbmenyn:  
Redigera förteckning  
Det här kommandot öppnar dialogrutan där du kan redigera förteckningen.  
Radera förteckning  
Med hjälp av det här kommandot raderar du den aktuella förteckningen.  
Alla förteckningar  
Då spelar det ingen som helst roll var markören befinner sig, i motsats till vad som gäller för kommandot Aktuell förteckning:  
Radnumrering  
Med den här funktionen kan du aktivera och konfigurera visningen av radnummer för ett dokument.  
Numrering på  
Om den här kryssrutan är markerad är radnumreringen aktiverad.  
Visa  
I det här området bestämmer du hur radnumreringen ska visas.  
Teckenformatmall  
Här kan du ställa in en teckenformatmall för numreringen.  
Du kan använda den eller välja en annan mall.  
I kombinationsfältet kan du välja bland samtliga tillgängliga teckenformatmallar, även de användardefinierade.  
Format  
Här kan du välja numreringsformat.  
Du kan välja mellan arabiska och romerska siffror eller bokstäver.  
Position  
Här placerar du radnumreringen i dokumentet.  
Med alternativen Till vänster och Till höger placerar du numreringen vid den vänstra eller högra kanten av textramen eller sidan.  
Effekten av alternativen Inre och Yttre beror på om det är raderna på en jämn eller udda sida i dokumentet som numreras.  
Avstånd  
Här ställer du in numreringens avstånd från styckeområdet eller textramen.  
Se till att inte ställa in för stort avstånd, för då riskerar du att inte se radnumren.  
Om du är osäker på hur mycket plats du har till förfogande, kan du orientera dig efter den horisontella linjalen ovanför arbetsområdet.  
Intervall...rader  
Här kan du ange i vilket intervall en radnumrering ska ske.  
Du kan t.ex. ange om varje, var femte eller var tionde rad ska numreras.  
Skiljetecken  
Förutom radnumret kan du definiera ett skiljetecken.  
Ett skiljetecken är ett valfritt tecken som visas mellan de numrerade raderna.  
Eftersom skiljetecken bara visas mellan radnumreringar, så är det meningslöst att ange ett skiljetecken om varje rad ska numreras.  
Text  
Här kan du skriva in ett valfritt tecken som ska visas som skiljetecken, t.ex. ett bindestreck ("-").  
Var...rad  
Här kan du ange skiljetecknets intervall.  
Om du t.ex. har lagt in en numrering för var tionde rad, kan du dessutom visa var femte rad med ett skiljetecken om du vill.  
Skiljetecken visas bara på sådana rader som saknar numrering.  
Om du ställer in samma värde här som du ställt in i området Visa under Intervall... rader har det ingen synlig effekt att ange ett skiljetecken.  
Räkna  
Här kan du ange om tomma rader och rader i textramar ska tas med i numreringen.  
Tomma rader  
Om du markerar den här rutan, räknas tomma rader vid radnumreringen.  
Rader i textram  
Markera den här rutan, om du även vill förse raderna i en textram med radnumrering.  
Numreringen av raderna i textramen sker oberoende av numreringen av raderna i dokumentet, och numreringen börjar med 1 i varje textram i dokumentet.  
Men när det gäller länkade ramar startar inte numreringen om i varje ram, utan löper oavbruten genom samtliga länkade ramar.  
Börja om på varje ny sida  
Markera den här rutan om numreringen ska börja om på varje sida.  
Uppdatera allt  
Med det här kommandot uppdaterar du hela dokumentet.  
Länkar, Fält, Alla förteckningar, Sidformatering.  
Fält  
Med det här kommandot uppdaterar du fältkommandon i det aktuella dokumentet.  
Länkar  
Med det här kommandot uppdaterar du länkarna i det aktuella dokumentet.  
När du har valt det här kommandot visas de uppdaterade versionerna av de länkade objekten i dokumentet.  
Alla diagram  
Med det här kommandot uppdaterar du alla diagram i dokumentet, vilkas tabelldata har ändrats.  
De uppdaterade diagrammen visas sedan i dokumentet.  
Uppdatera  
Här kan du bland annat genomföra en sidformatering manuellt samt uppdatera förteckningar.  
Numrering på / av  
Med den här ikonen tilldelar du de markerade styckena en numrering.  
För redan numrerade stycken upphävs numreringen när du klickar på ikonen.  
Med hjälp av objektlisten för numreringar kan du lätt och snabbt strukturera alla stycken.  
Du aktiverar numreringsobjektlisten med hjälp av pilknappen i den högra kanten av textobjektlisten.  
I onlinelayout är några av alternativen för numrering / punktuppställning inte tillgängliga.  
Numrering på / av  
Länka  
Med den här ikonen kan du länka ihop den markerade ramen med en annan efterföljande ram.  
Textinnehållet i länkade ramar bryts automatiskt från ram till ram.  
Länka  
Lös upp länkning  
Med den här ikonen upphäver du länkningen av en ram till dess efterföljare.  
Du kan välja att enbart bryta kedjan till efterföljaren och inte till föregångaren.  
Därför kan du bara aktivera ikonen Lös upp länkning om du har markerat en länkad föregångar-ram.  
Lös upp länkning  
Infoga rad  
När du klickar på den här ikonen, infogar du exakt en rad i tabellen nedanför markörens position.  
Du kan infoga flera rader samtidigt om du öppnar dialogrutan Infoga rader via menykommandot Format - Rad - Infoga, eller om du markerar flera rader innan du klickar på ikonen.  
I det sistnämnda fallet får de infogade raderna samma relativa höjder som de markerade raderna.  
Infoga rad  
Infoga kolumn  
När du klickar på den här ikonen, infogar du en kolumn i tabellen efter markörens position.  
Du kan infoga flera kolumner samtidigt om du öppnar dialogrutan via menykommandot Format - Kolumn - Infoga..., eller om du markerar flera kolumner innan du klickar på ikonen.  
I det senare fallet får de infogade kolumnerna samma relativa bredder som de markerade kolumnerna.  
Infoga kolumn  
Optimera  
Med den här ikonen öppnar du en utrullningslist med olika funktioner för optimering av tabellrader och -kolumner.  
Ikon på objektlisten:  
Optimera  
Du kan välja följande funktioner:  
Optimal radhöjd  
Optimal kolumnbredd  
Tabell: fast  
Om det här läget är aktivt och du ändrar en rad och / eller kolumn, så påverkar detta bara den intilliggande raden / kolumnen.  
Tabell: fast  
Tabell: fast, proportionell  
Om det här läget är aktivt och du ändrar en rad och / eller kolumn, så påverkar det hela tabellen.  
Tabell: fast, proportionell  
Tabell: variabel  
Om det här läget är aktivt och du ändrar en rad och / eller kolumn, så påverkar det tabellstorleken.  
Tabell: variabel  
Summa  
När du klickar på den här ikonen på tabellobjektlisten startar du summafunktionen.  
Sätt först cellmarkören i cellen eller markera cellerna där summaformeln ska föras in.  
Om cellerna redan är fyllda med data, registrerar %PRODUCTNAME mestadels automatiskt för vilket cellområde du vill använda summafunktionen.  
Klicka på ikonen Överta om du vill överta summaformeln så som den visas på inmatningsraden.  
Den här ikonen visas bara om du inte har aktiverat inmatningsraden.  
Summa  
Numrering av  
Med den här ikonen tar du bort automatisk numrering / punktuppställning i det aktuella stycket eller i de markerade styckena.  
Numrering av  
Nedåt med undernivåer  
Med den här ikonen flyttar du styckena tillsammans med alla underordnade stycken en nivå nedåt.  
Den visas bara om markören står i en punktuppställning eller numrering.  
Nedåt med undernivåer  
Uppåt med undernivåer  
Med den här ikonen flyttar du styckena tillsammans med alla underordnade stycken en nivå uppåt.  
Den visas bara om markören står i en punktuppställning eller numrering.  
Uppåt med undernivåer  
Infoga post utan nummer  
Med hjälp av den här ikonen kan du infoga ett stycke utan numrering på den aktuella nivån.  
Den befintliga numreringen påverkas inte.  
Ikonen visas bara om markören står i en punktuppställning eller numrering.  
Infoga post utan nummer  
Flytta uppåt med undernivåer  
Med den här ikonen placerar du ett stycke med alla understycken framför föregående stycke.  
Den visas bara om markören står i en punktuppställning eller numrering.  
Flytta uppåt med undernivåer  
Flytta nedåt med undernivåer  
Med den här ikonen placerar du ett stycke med alla underordnade stycken efter följande stycke.  
Den visas bara om markören står i en punktuppställning eller numrering.  
Flytta nedåt med undernivåer  
Starta om numrering  
Den här ikonen startar om en numrering.  
Den visas bara om markören står i en punktuppställning eller numrering.  
Starta om numrering  
Sidnummer  
I det här fältet på statuslisten visas aktuellt sidnummer.  
Om du dubbelklickar på fältet öppnas Navigator med vars hjälp du kan navigera i dokumentet.  
Om du högerklickar visas alla bokmärken i dokumentet.  
Du kan klicka på ett om du vill placera markören där.  
Den visade sidan (x) och det totala antalet sidor (y) i dokumentet visas i form av Sida x / y.  
Om du bläddrar med musen genom ett flersidigt dokument visas här numret på den sida som visas när du släpper musknappen.  
Om du flyttar knappen på den högra bildrullningslisten visas sidnumren som tipshjälp.  
Formateringen av sidnumreringen på statuslisten och bildrullningslisten är identisk och så som du har definierat den.  
Om du dubbelklickar på det här fältet visas eller döljs Navigator.  
Om du vill gå till en viss sida med hjälp av Navigator, anger du sidnumret i rotationsfältet Sida i Navigator och trycker på Retur.  
Med tangentkombinationen Skift + Kommando Ctrl +F5 växlar du till inmatning av sidnummer.  
När du trycker på Retur, flyttas visning och markör till början av den valda sidan.  
Kombinerad visning  
I det här fältet visas aktuella upplysningar om dokumentet.  
Om textmarkören exempelvis står i ett namngivet område, visas namnet på området här.  
Om markören står i en tabell, visas namnet på tabellcellen.  
När du redigerar ramar eller ritelement visas objektets storlek här.  
Här kan du ange ett fältkommando, som infogas i dokumentet där markören står för tillfället.  
Om markören står i en tabell öppnar du dialogrutan Tabellformat genom att dubbelklicka i det här fältet.  
På motsvarande sätt kan du här, beroende på vilket objekt som är markerat, öppna en dialogruta för att redigera ett område, ett grafikobjekt, en ram, ett OLE-objekt, en direkt numrering eller ritobjekts position och storlek.  
Utföra eller redigera hyperlänkar  
I det här fältet på statuslisten växlar du mellan Utför (HYP) och Redigera (SEL) för text-hyperlänkarna i dokumentet genom att klicka med musen.  
Visning:  
Verkan:  
HYP  
Om du klickar på en hyperlänk laddas den URL som den innehåller.  
SEL  
Du kan klicka på en hyperlänktext som på normal text och redigera den.  
Om Du inte vill redigera den synliga texten i hyperlänken, utan URL:en, så måste HYP visas i detta fält på statuslisten.  
Då kan du peka på hyperlänken, trycka på musknappen och hålla ner den medan du drar till hyperlänklisten.  
Där kan du redigera både text och länk (URL).  
Med knappen Länk infogar du den redigerade hyperlänken vid textmarkörens position i dokumentet.  
Om Du inte har infogat hyperlänken som text, utan som kommandoknapp (se knappen Länk), så kan Du redigera hyperlänken enbart genom att ändra kontrollfältets egenskaper:  
Markera kommandoknappen och anropa kommandot Kontrollfält... via snabbmenyn.  
I kommandoknappens Egenskapsdialogruta kan Du både redigera den synliga texten på knappen och URL:en.  
Förhandsgranskning: två sidor  
Om du klickar på den här ikonen visas två sidor i förhandsgranskningsfönstret.  
Udda numrerade sidor står alltid till höger, jämna till vänster.  
Förhandsgranskning: två sidor  
Förhandsgranskning: fyra sidor  
Om du klickar på den här ikonen visas fyra sidor i fönstret för förhandsgranskning.  
Förhandsgranskning: fyra sidor  
Skala  
Klicka på den här ikonen om du vill ändra antalet sidor som visas på bildskärmen.  
Om du klickar snabbt på den öppnas en dialogruta, där du kan bestämma hur de olika sidorna ska visas vid förhandsgranskningen.  
De inställningar som Du gör i dialogrutan kan Du på ett enkelt sätt även göra med hjälp av musen:  
Då öppnas en popup-listruta, där Du kan ange det antal sidor som ska visas med musen.  
Gå med musen över önskat antal rader och kolumner (en rad och en kolumn motsvarar en sida) och bekräfta Ditt val genom att klicka med musen.  
Skala  
Visa  
I dialogrutan visas två rotationsfält, där Du kan ange det antal sidor som ska visas.  
Vid en rad och en kolumn visas exakt en sida, vid en rad och två kolumner visas en dubbelsida, dvs vänster och höger sida tillsammans.  
Rader  
Här ställer Du in antalet rader av sidor under varandra.  
Kolumner  
Här ställer Du in antalet kolumner av sidor bredvid varandra.  
Skriv ut förhandsgranskning  
Om du klickar på den här ikonen skrivs förhandsgranskningen ut.  
Förhandsgranskningen skrivs ut i den form som visas på bildskärmen.  
Tillsammans med menyn Visa - Skala kan du här ange att du skriver ut förhandsvisningar med t.ex. 8 sidor bredvid varandra och 10 sidor under varandra av ett flersidigt dokument, om du vill få en överblick över uppdelningen av text till grafik eller liknande.  
Skriv ut förhandsgranskning  
Utskriftsalternativ förhandsgranskning  
Om du klickar på den här ikonen öppnas en dialog där du kan göra inställningar för utskriften av dina dokumentsidor.  
Du kan också öppna dialogen via snabbmenyn (här heter kommandot Skrivaralternativ).  
Sidorna förminskas jämnt vilket kan leda till att inte hela arket utnyttjas vid utskriften och en kant lämnas kvar om det är ett textdokument på flera sidor.  
Inställningarna som Du har gjort i dialogrutan Utskriftsalternativ gäller bara om dokumentet skrivs ut via kommandoknappen Skriv ut förhandsgranskning.  
Utskriftsalternativ förhandsgranskning  
Uppdelning  
I det här området ställer Du in resp. anger antalet rader och kolumner som ska skrivas ut.  
Om flera dokumentsidor ska skrivas ut på en sida bestämmer Du antalet dokumentsidor som ska ligga över och bredvid varandra.  
Även om Ditt dokument bara består av en sida, kan Du bestämma storleken på utskriften här.  
Rader  
Med de här rotationsknapparna definierar Du antalet rader, d.v.s. dokumentsidorna som ligger över varandra.  
Kolumner  
Med de här rotationsknapparna bestämmer Du antalet kolumner, d.v.s. dokumentsidor som ligger bredvid varandra.  
Marginaler  
I det här området bestämmer Du marginalerna på utskriftssidan.  
Vänster  
Du betsämmer hur bred den vänstra marginalen ska vara med rotationsknapparna.  
Uppåt  
Du bestämmer hur bred den övre marginalen ska vara med rotationsknapparna.  
Höger  
Du bestämmer hur bred den högra marginalen ska vara med rotationsknapparna.  
Nedåt  
Du bestämmer hur bred den undre marginalen ska vara med rotationsknapparna.  
Avstånd  
I området avstånd definierar Du de horisontella och vertikala avstånden mellan de förminskade dokumentsidorna på utskriftssidan.  
Horisontell  
Använd de här rotationsknapparna till att definiera ett vågrätt avstånd.  
Vertikalt  
Använd de här rotationsknapparna till att definiera ett lodrätt avstånd.  
Format  
I det här området bestämmer Du vilket format utskriften ska ha.  
Liggande  
Välj det här alternativfältet om Du vill skriva ut i liggande format.  
Stående  
Välj det här alternativfältet om Du vill skriva ut i stående format.  
Standard  
Om Du klickar på den här kommandoknappen används inte något fast antal rader och kolumner för utskriften av förhandsgranskningen, utan det antal som för tillfället visas i förhandsgranskningen.  
Cellreferens  
I det här fältet visas cellmarkörens position i en tabell.  
Cellreferens  
Formel  
Från undermenyn till den här ikonen kan du infoga en formel.  
Sätt markören i tabellen i cellen eller i dokumentet på det ställe där resultatet ska visas.  
Klicka sedan på den här ikonen, och välj önskad formel från undermenyn.  
Formeln infogas på inmatningsraden.  
Om du vill välja ett område med celler i en textdokumenttabell markerar du cellerna i tabellen.  
Korrekt cellreferens infogas på inmatningsraden.  
Infoga fler parametrar som behövs och avsluta inmatningen genom att klicka på ikonen Överta.  
Naturligtvis kan du också mata in formeln direkt, så snart du känner till syntaxen (det är till exempel nödvändigt i dialogrutornas inmatningsfält för Fältkommandon och Redigera fältkommando).  
Ikon på formellisten:  
Formel-undermeny  
Formelelementens tabeller  
De fyra räknesätten  
Addition  
+  
Beräknar summan.  
Exempel: <A1> + 8  
Subtraktion  
-  
Beräknar differensen.  
Exempel:  
10 - <B5>  
Multiplikation  
MUL eller *  
Beräknar produkten.  
Exempel:  
7 MUL 9  
Division  
DIV eller /  
Beräknar kvoten.  
Exempel:  
100 DIV 1,15  
Grundfunktioner på undermenyn  
Summa  
SUM  
Beräknar summan av de markerade cellerna.  
Exempel:  
SUM <A2:C2> visar summan av värdena i cellerna från A2 till C2  
Avrunda  
ROUND  
Avrundar ett tal till ett angivet antal decimaler.  
Exempel:  
15,678 ROUND 2 visar 15,68  
Procent  
PHD  
Beräknar ett procentvärde.  
Exempel:  
10 + 15 PHD visar 11,50  
Kvadratrot  
SQRT  
Beräknar kvadratroten.  
Exempel:  
SQRT 25 visar 5,00  
Upphöja  
POW  
Beräknar potensen.  
Exempel:  
2 POW 8 visar 256,00  
Operatorer  
Här kan du använda operatorer.  
Operatorer  
Listavgränsare  
_BAR_  
Skiljer elementen i listor från varandra.  
Exempel på en lista:  
10_BAR_ 20_BAR_50_BAR_<C6>_BAR_<A2:B6> _BAR_20  
Lika med  
EQ eller ==  
Testar likhet.  
Om inte lika med, är resultatet 0 (falskt), annars 1 (sant).  
Exempel: <A1> EQ 2 visar 1, om innehållet i A1 är lika med 2.  
Inte lika med  
NEQ eller !=  
Testar olikhet.  
Exempel: <A1> NEQ 2 visar 0 (falskt), om innehållet i A1 är lika med 2.  
Mindre än eller lika med  
LEQ  
Testar mindre än eller lika med.  
Exempel: <A1> LEQ 2 visar 1 (sant), om innehållet i A1 är mindre än eller lika med 2.  
Större än eller lika med  
GEQ  
Testar större än eller lika med.  
Exempel: <A1> GEQ 2 visar 1 (sant), om innehållet i A1 är större eller lika med 2.  
Mindre än  
L  
Testar mindre än.  
Exempel: <A1> L 2 visar 1 (sant), om innehållet i A1 är mindre än 2.  
Större än  
G  
Testar större än.  
Exempel: <A1> G 2 visar 1 (sant), om innehållet i A1 är större än 2.  
Logiskt Eller  
OR  
Testar logiskt Eller.  
Exempel:  
0 OR 0 visar 0 (falskt), allt annat visar 1 (sant)  
Logiskt Exklusivt Eller  
XOR  
Testar logiskt Exklusivt Eller.  
Exempel:  
1 XOR 0 visar 1 (sant)  
Logiskt Och  
AND  
Testar logiskt Och.  
Exempel:  
1 AND 2 visar 1 (sant)  
Logiskt Inte  
NOT  
Testar logiskt Inte.  
Exempel:  
NOT 1 (sant) visar 0 (falskt)  
Statistiska funktioner  
Några enkla statistiska funktioner står till förfogande.  
Medelvärde  
MEAN  
Beräknar det aritmetiska medelvärdet i ett område eller en lista.  
Exempel:  
MEAN 10_BAR_ 30 _BAR_20 visar 20,00  
Minimum  
MIN  
Beräknar det minsta värdet i en lista eller ett område.  
Exempel:  
MIN 10_BAR_ 30 _BAR_20 visar 10,00  
Maximum  
MAX  
Beräknar det största värdet i en lista eller ett område.  
Exempel:  
MAX 10_BAR_ 30 _BAR_20 visar 30,00  
Trigonometriska funktioner  
Här kan du välja mellan trigonometriska funktioner.  
sinus  
SIN  
Beräknar sinus i radianer.  
Exempel:  
SIN (PI / 2)  
cosinus  
COS  
Beräknar cosinus i radianer.  
Exempel:  
COS 1  
tangens  
TAN  
Beräknar tangens i radianer.  
Exempel:  
TAN <A1>  
arcussinus  
ASIN  
Beräknar arcussinus i radianer.  
Exempel:  
ASIN 1  
arcuscosinus  
ACOS  
Beräknar arcuscosinus i radianer.  
Exempel:  
ACOS 1  
arcustangens  
ATAN  
Beräknar arcustangensen i radianer.  
Exempel:ATAN 1  
Variabler för dokumentegenskaper  
De följande egenskaperna för ett dokument finns även under Arkiv - Egenskaper - Statistik.  
CHAR  
Antal tecken i dokumentet  
WORD  
Antal ord i dokumentet  
PARA  
Antal stycken i dokumentet  
GRAF  
Antal grafikobjekt i dokumentet  
TABLES  
Antal tabeller i dokumentet  
OLE  
Antal OLE-objekt i dokumentet  
PAGE  
Totalt antal sidor i dokumentet  
Andra definierade värden  
Pi  
PI  
3,1415...  
Eulers tal  
E  
2,7182...  
Sant  
TRUE  
inte lika med 0  
Falskt  
FALSE  
0  
Avbryt  
Om du klickar på den här ikonen tas innehållet i inmatningsraden bort och formellisten stängs.  
Avbryt  
Överta  
Genom att klicka på den här ikonen övertar du innehållet på inmatningsraden och stänger formellisten.  
Innehållet på inmatningsraden infogas vid markörens position i dokumentet.  
Överta  
Formelområde  
I den här delen av formellisten bygger du upp formeln, antingen genom att skriva in formeln direkt eller genom att ta formelikonens popupmeny till hjälp.  
Formelområde  
Infoga  
Om du klickar något längre öppnas en utrullningslist med olika funktioner för infogning av ramar, grafikobjekt, tabeller o.s.v.  
Om du klickar kort aktiveras verktyget som visas som ikon.  
Ikon på verktygslisten:  
Infoga  
När du har valt en funktion på utrullningslisten för första gången, visas alltid ikonen för den senast infogade funktionen på verktygslisten.  
Du kan välja följande funktioner:  
Infoga ram manuellt  
Infoga grafik  
Infoga tabell  
Dokument  
Infoga fotnot direkt  
Infoga slutnot direkt  
Infoga specialtecken  
Infoga område  
Infoga indexmarkering  
Infoga bokmärke  
Infoga fältkommandon (HTML-dokument)  
Med den här ikonen öppnar du en undermeny där du kan infoga fältkommandon.  
Håll ner musknappen lite längre på ikonen och välj önskat fältkommando.  
Om du klickar kort öppnas dialogrutan Fältkommandon.  
Du kan välja följande funktioner:  
Andra...  
Datum  
Här infogar du aktuellt datum som fältkommando.  
Datumet uppdateras inte automatiskt.  
Om du vill ha ett annat datumformat eller en automatisk anpassning av datumet, väljer du kommandot Infoga - Fältkommando - Andra... för att infoga fältkommandot och gör önskade inställningar i dialogrutan Fältkommandon.  
Men du kan också ändra formatet för ett redan infogat datumfält med hjälp av menykommandot Redigera - Fältkommando....  
Klockslag  
Här infogar du aktuellt klockslag som fältkommando.  
Det hämtas från operativsystemets systeminställningar.  
För formatering används ett standardformat.  
Du kan inte anpassa tidsangivelsen genom att uppdatera fältkommandot med F9.  
Om du vill ha ett annat tidsformat eller möjlighet att anpassa klockslaget, väljer du kommandot Infoga - Fältkommando - Andra... för att infoga fältkommandot och gör önskade inställningar i dialogrutan Fältkommandon.  
Men du kan också ändra formatet för ett redan infogat klockslagsfält med hjälp av menykommandot Redigera - Fältkommando....  
Sidnummer  
Här infogar du aktuellt sidnummer som fältkommando vid markörens position.  
Standardformatet hämtas från sidformatmallen.  
Om du vill ha ett annat format eller möjlighet att korrigera sidnumret, väljer du kommandot Infoga - Fältkommando - Andra... för att infoga fältkommandot och gör önskade inställningar i dialogrutan Fältkommandon.  
Men du kan också ändra formateringen och korrigeringsvärdet i fältet som du har infogat med menykommandot Sidnummer med hjälp av menykommandot Redigera - Fältkommando....  
Sidantal  
Här infogar du dokumentets totala antal sidor som fältkommando.  
För detta används standardmässigt arabiska siffror.  
Om du vill ha ett annat visningsformat för sidantalet, väljer du kommandot Infoga - Fältkommando - Andra... för att infoga fältkommandot och gör önskade inställningar i dialogrutan Fältkommandon.  
Men du kan även ändra formateringen i fältet som du infogat med menykommandot Sidantal med hjälp av menykommandot Redigera - Fältkommando....  
Ämne  
Här infogar du det som dokumentegenskap angivna ämnet som fältkommando.  
Fältkommandot övertar då posten som finns under Arkiv - Egenskaper - Beskrivning i fältet Ämne.  
Om du vill infoga en annan dokumentegenskap som fältkommando, väljer du kommandot Infoga - Fältkommando - Andra... och gör önskade inställningar i dialogrutan Fältkommandon.  
Här hittar du samtliga tillgängliga fälttyper under fliken Dokumentinfo.  
Rubrik  
Här infogar du den som dokumentegenskap angivna rubrik som fältkommando.  
Fältkommandot övertar då den post som du sparat under Arkiv - Egenskaper - Beskrivning i fältet Rubrik.  
Om du vill infoga en annan dokumentegenskap som fältkommando, väljer du kommandot Infoga - Fältkommando - Andra... och gör önskade inställningar i dialogrutan Fältkommandon.  
Du hittar samtliga tillgängliga fälttyper under fliken Dokumentinfo.  
Författare  
Här infogar du användarnamnet som fältkommando.  
Fältkommandot övertar då den post som finns under Verktyg - Alternativ - %PRODUCTNAME - Användardata.  
Grafik  
Bara tomma ramar visas som platshållare.  
Grafik  
Direktmarkör på / av  
Med den här ikonen sätter du på eller stänger av direktmarkören.  
Med direktmarkören kan du klicka på ett valfritt ställe i dokumentet och börja skriva där.  
Om du öppnar dialogrutan för direktmarkörens egenskaper under Verktyg - Alternativ - Textdokument - Markör, kan du ange hur texten infogas vid den position där du klickar.  
Direktmarkör på / av  
Med direktmarkören kan du, förutom att placera text på en valfri position i dokumentet, bestämma infogningspositionen för grafiska objekt, tabeller, ramar och andra objekt genom att klicka med musen.  
Om du placerar direktmarkören ungefär i mitten mellan den vänstra och högra kanten på en sida eller tabellcell, så centreras den infogade texten.  
På motsvarande sätt kan du mata in den följande texten högerjusterat när du har placerat direktmarkören vid den högra kanten.  
När du har aktiverat AutoKorrigering och infogar tomma stycken, tabbar och blanksteg med direktmarkören, kan det hända att de direkt tas bort automatiskt.  
De kan nämligen inte användas samtidigt.  
Direktmarkören placerar markören med hjälp av tabbar.  
Om du ändrar tabbarna i efterhand, t.ex. genom att tilldela en annan styckeformatmall, så kan detta ändra textens position på sidan.  
Infoga sidhuvud  
Om du klickar på den här ikonen infogar du ett sidhuvud i HTML-dokumentet.  
Infoga sidhuvud  
Infoga sidfot  
Om du klickar på den här ikonen infogar du en sidfot i HTML-dokumentet.  
Infoga sidfot  
Infoga  
Om du håller ner musknappen öppnas en utrullningslist med olika funktioner för infogning av grafiska objekt, tabeller, dokument, specialtecken o.s.v.  
Om du klickar snabbt, aktiveras det verktyg som visas som ikon.  
Ikon på verktygslisten:  
Infoga  
När du har valt en funktion på utrullningslisten för första gången, visas ikonen för den senast infogade funktionen på verktygslisten.  
Du kan välja följande funktioner:  
Infoga ram manuellt  
Grafik  
Tabell  
Dokument  
Specialtecken  
Infoga område  
Bokmärke  
Infoga fältkommandon  
Med den här ikonen öppnar du en undermeny där du kan infoga viktiga fältkommandon.  
Håll ner musknappen på ikonen och välj det önskade fältkommandot.  
Om du klickar snabbt, öppnas dialogrutan Fältkommandon.  
Ikon på verktygslisten:  
Du kan välja följande funktioner:  
Andra...  
Animerad text  
Animerad text  
Kortkommandon för textdokument  
Här hittar du en förteckning över tangentkombinationer som du har användning för i textdokument.  
Dessutom gäller de allmänna tangentkombinationerna i %PRODUCTNAME.  
Funktioner i textdokument med funktionstangenterna  
Tangentkombination  
Effekt  
F2  
Formellist  
Kommando Ctrl +F2  
Infoga fältkommando  
F3  
Expandera AutoText  
Kommando Ctrl +F3  
Redigera AutoText  
F4  
Öppna datakällvy  
F5  
Navigator på / av  
Skift+F5  
Hoppa till nästa ram  
Kommando Ctrl +Skift+F5  
Aktivera Navigator  
F7  
Rättstavningskontroll  
Kommando Ctrl +F7  
Synonymordlista  
F8  
Utvidgningsläge  
Kommando Ctrl +F8  
Markeringar på / av  
Skift+F8  
Kompletteringsläge  
F9  
Uppdatera fält  
Kommando Ctrl +F9  
Visa fältkommandon  
Skift+F9  
Beräkna tabell  
Kommando Ctrl +Skift+F9  
Uppdatera inmatningsfält  
Kommando Ctrl +F10  
Kontrolltecken på / av  
F11  
Stylist på / av  
Skift+F11  
Skapa formatmall  
Kommando Ctrl +Skift+F11  
Uppdatera formatmall  
F12  
Numrering på  
Kommando Ctrl +F12  
Infoga tabell  
Skift+F12  
Punktuppställning på  
Kommando Ctrl +Skift+F12  
Numrering / punktuppställning av  
Speciella tangentstyrningar för textdokument  
Tangentkombination  
Effekt  
Kommando Ctrl +A  
Markera allt  
Kommando Ctrl +B  
Marginaljustering  
Kommando Ctrl +D  
Dubbel understrykning  
Kommando Ctrl +E  
Centrerad  
Kommando Ctrl +G  
Sök och ersätt  
Kommando Ctrl +H  
Upphöjd  
Kommando Ctrl +L  
Vänsterjusterad  
Kommando Ctrl +R  
Högerjusterad  
Kommando Ctrl +T  
Nedsänkt  
Kommando Ctrl +Y  
Mallkatalog  
Kommando Ctrl +1  
Enkelt radavstånd  
Kommando Ctrl +2  
Dubbelt radavstånd  
Kommando Ctrl +5  
1,5 radavstånd  
Kommando Ctrl +  
Beräknar det markerade området (t.ex. 3487+3456).  
Resultatet kopieras till urklippet och måste klistras in därifrån.  
Kommando Ctrl -  
Användardefinierat bindestreck; ett bindestreck som du har infogat i ordet.  
Kommando Ctrl +Skift -  
Skyddat bindestreck (används inte som bindestreck vid avstavning)  
Kommando Ctrl * (bara tecken på den numeriska delen av tangentbordet)  
Utföra makrofält  
Kommando Ctrl +mellanslag  
Fast mellanrum.  
Fasta mellanrum bryts inte i slutet av raden och marginaljusteras inte.  
Skift+Retur  
Radbrytning utan nytt stycke  
Kommando Ctrl +Retur  
Manuell sidbrytning  
Kommando Ctrl +Skift+Retur  
Kolumnbrytning i texter med flera kolumner  
Alternativ Alt +Retur  
Infogar nytt stycke utan punktuppställningstecken i punktuppställning  
Alternativ Alt +Retur  
Infogar ett stycke direkt före eller efter ett område  
Vänsterpil  
Insättningspunkten åt vänster  
Skift+Vänster piltangent  
Insättningspunkten åt vänster med markering  
Kommando Ctrl +Vänster piltangent  
Hoppa till ordets början  
Kommando Ctrl +Skift+Vänster piltangent  
Markera ord för ord åt vänster  
Högerpil  
Insättningspunkten åt höger  
Skift+Höger piltangent  
Insättningspunkten åt höger med markering  
Kommando Ctrl +Höger piltangent  
Hopp till ordets slut  
Kommando Ctrl +Skift+Höger piltangent  
Markera ord för ord åt höger  
Övre piltangent  
Rad uppåt  
Skift+Övre piltangent  
Rad uppåt med markering  
Nedre piltangent  
Rad nedåt  
Skift+Nedre piltangent  
Rad nedåt med markering  
Home  
Hopp till början av raden  
Skift+Home  
Hopp till början av raden med markering  
End  
Hopp till slutet av raden  
Skift+End  
Hopp till slutet av raden med markering  
Kommando Ctrl +Home  
Hopp till början av dokumentet  
Kommando Ctrl +Skift+Home  
Hopp till början av dokumentet med markering  
Kommando Ctrl +End  
Hopp till slutet av dokumentet  
Kommando Ctrl +Skift+End  
Hopp till slutet av dokumentet med markering  
Kommando Ctrl +PageUp  
Flytta markören mellan text och sidhuvud  
Kommando Ctrl +PageDown  
Flytta markören mellan text och sidfot  
Insert  
Infogningsläge på / av  
PageUp  
Bildskärmssida uppåt  
Skift+PageUp  
Bildskärmssida uppåt med markering  
PageDown  
Bildskärmssida nedåt  
Skift+PageDown  
Bildskärmssida nedåt med markering  
Kommando Ctrl +Delete  
Raderar text till ordets slut  
Kommando Ctrl +Backsteg  
Raderar text till ordets början  
Kommando Ctrl +Skift+Delete  
Raderar text till meningens slut  
Kommando Ctrl +Skift+Backsteg  
Raderar text till meningens början  
Kommando Ctrl +Tabb  
Vid automatisk ordkomplettering: nästa förslag  
Kommando Ctrl +Skift+Tabb  
Vid automatisk ordkomplettering: föregående förslag  
Alternativ Alt +O  
I dialogrutan Rättstavning:  
Det ord som ursprungligen har markerats som okänt / felaktigt (Original) övertas på inmatningsraden (Ord)  
Kommando Ctrl +Dubbelklick med musen  
Använd denna kombination om du snabbt vill förankra eller frigöra Navigator, Stylist eller andra fönster.  
Flytta stycken och överskrifter  
Numreringar anpassas automatiskt  
Tangentkombination  
Effekt  
Kommando Ctrl +Övre piltangent  
Flytta aktuellt stycke eller markerade stycken ett stycke uppåt.  
Kommando Ctrl +Nedre piltangent  
Flytta aktuellt stycke eller markerade stycken ett stycke nedåt.  
Tabb  
Överskriften i formatet "Överskrift X" (X = 1-9) flyttas ned en nivå i dispositionen.  
Skift+Tabb  
Överskriften i formatet "Överskrift X" (X = 2-10) flyttas upp en nivå i dispositionen.  
Kommando Ctrl +Tabb  
I början av en överskrift: infogar en tabb.  
För att du ska kunna växla överskriftsnivåer med hjälp av tangentbordet, måste du placera markören framför överskriften innan du trycker på tangenterna.  
Kortkommandon i tabeller  
Tangentkombination  
Effekt  
Kommando Ctrl +A  
Om den aktuella cellen är tom:  
Markerar hela tabellen.  
Annars:  
Markerar innehållet i den aktuella cellen, en förnyad aktivering markerar hela tabellen  
Kommando Ctrl +Home  
Om den aktuella cellen är tom:  
Hoppar till början av tabellen.  
Annars:  
Hoppar vid första tryckningen till början av den aktuella cellen, vid nästa tryckning till början av den aktuella tabellen, vid tredje tryckningen till början av dokumentet.  
Kommando Ctrl +End  
Om den aktuella cellen är tom:  
Hoppar till slutet av tabellen.  
Annars:  
Hoppar vid första tryckningen till slutet av den aktuella cellen, vid nästa tryckning till slutet av den aktuella tabellen, vid tredje tryckningen till slutet av dokumentet.  
Kommando Ctrl +Tabb  
Infogar en tabb (bara i tabeller)  
Kommando Ctrl +Skift+Övre piltangent  
Början av tabellen  
Kommando Ctrl +Skift+Nedre piltangent  
Slutet av tabellen  
Alternativ Alt +Piltangent  
Förstorar / förminskar kolumnen / raden vid högra / nedre cellkanten  
Alternativ Alt +Skift+Piltangent  
Förstorar / förminskar kolumnen / raden vid vänstra / övre cellkanten  
Alternativ+Kommando Alt+Ctrl +Piltangent  
Som Alternativ Alt, bara den aktuella cellen förändras  
Alternativ+Kommando Alt+Ctrl +Skift+Piltangent  
Som Alternativ Alt, bara den aktuella cellen förändras  
Alternativ Alt +Insert  
3 sekunder i infogningsläge, piltangenten infogar rad / kolumn, Kommando Ctrl +piltangent infogar cell  
Alternativ Alt +Delete  
3 sekunder i raderingsläge, piltangenten raderar rad / kolumn, Kommando Ctrl +piltangent sammanfogar cell med granncell till en cell  
Kommando Ctrl +Skift+T  
Upphäver cellskyddet i alla markerade tabeller.  
Om markören står någonstans i dokumentet, d.v.s. om ingen tabell har markerats, upphävs cellskyddet för alla tabeller.  
Skift Kommando +Ctrl +Delete  
Om du inte har markerat något, raderas nästa cellinnehåll.  
Om du har markerat celler, raderas hela raderna inom markeringen.  
Om du har markerat samtliga rader helt eller delvis, raderas hela tabellen.  
Flyttning och storleksändring av ramar / grafikobjekt och objekt  
Tangentkombination  
Effekt  
Alternativ Alt +Piltangent  
Flytta objekt.  
Alternativ+Kommando Alt+Ctrl +Piltangent  
Storleksändring genom att den högra / nedre kanten flyttas.  
Alternativ+Kommando Alt+Ctrl +Skift+Piltangent  
Storleksändring genom att den vänstra / övre kanten flyttas.  
Placera objekt  
Objekten på en textsida, som t.ex. grafikobjekt och textramar, kan du förankra på olika sätt.  
Här presenteras de olika möjligheterna med en ram som exempel:  
Förankring  
Effekt  
som tecken  
Ramen står som ett tecken i texten och påverkar alltså radhöjd och brytning.  
vid tecken  
Ramen är fast knuten till ett tecken med sina X - och Y-koordinater, t.ex. alltid vid sidmarginalen i X-riktningen och alltid på tecknets höjd i y-riktningen (Marginalram).  
Ramen ska ha inställningen "Genomflöde".  
vid stycke  
Ramen är fast knuten till ett stycke och placeringen rättas efter stycket.  
vid sida  
Ramen har alltid samma placering i förhållande till sidmarginalerna.  
vid ram  
Ramen har en fast placering innanför den överordnade ramen.  
Det går också att välja placeringen i förhållande till förankringen med olika alternativ.  
Det är t.ex. möjligt att sätta ramen vid en fast position i förhållande till sidmarginalen, styckemarginalen, textområdet och så vidare.  
Rampositionen kan spegelvändas automatiskt på jämna sidor så att en fast position i förhållande till den högra sidmarginalen blir en spegelvänd position vid den vänstra sidmarginalen.  
På det här sättet kan du t.ex. alltid placera ett grafikobjekt vid den inre kanten av sidans yttre marginal.  
Om grafikobjektet t.ex. är en pil som pekar på texten, är det praktiskt att spegelvända den automatiskt på jämna sidor.  
Då använder du alternativet spegelvänd på jämna sidor under fliken Typ i dialogrutan Grafik (meny Format - Grafik).  
Kapitel i Navigator  
Här kan du ändra ordningen på kapitel eller deras nivå i hierarkin av kapitel och underordnade kapitel.  
Det enda villkoret för att detta ska fungera är att du har försett kapitelrubrikerna med styckeformatmallarna för överskrifter (eller ange de styckeformatmallar som du har valt för överskrifterna under Verktyg - Kapitelnumrering).  
Navigator som fritt fönster eller förankrat  
Håll ner Kommando Ctrl -tangenten och dubbelklicka på det gråa området i kanten av Navigator, t.ex. bredvid eller under ikonerna.  
Navigator förankras i fönsterkanten eller blir till ett fritt fönster igen, vars storlek och placering du kan bestämma genom att dra med musen.  
Placering och storlek registreras automatiskt.  
Du växlar mellan förankrat och fritt Navigatorfönster genom att dubbelklicka.  
Om du dubbelklickar på en överskrift i Navigator placeras textmarkören på motsvarande ställe i texten.  
Du kan ändra placeringen av kapitel med dra-och-släpp.  
Du kan också använda ikonerna Kapitel uppåt och Kapitel nedåt.  
Kapitlens innehåll och deras underordnade kapitel flyttas naturligtvis också.  
Om du håller ner Kommando Ctrl -tangenten när du drar och släpper kan du flytta kapitelöverskrifterna utan deras innehåll. (Ikonen Draläge påverkar bara dra-och-släpp mellan Navigator och dokument).  
Du ställer in detta med ikonen Visade överskriftsnivåer i Navigator.  
AutoText med AutoComplete  
1.  
Markera rutan Visa resten av namnet som tips vid inmatningen i dialogrutan AutoText.  
2.  
Från och med den tredje likadana bokstaven visas en tipshjälp med hela namnet från AutoText.  
3.  
Du infogar AutoText-blocket genom att trycka på Retur.  
Om det finns flera AutoText-namn som börjar likadant i tipshjälpen kan du bläddra framåt bland AutoText-namnen med Kommando Ctrl +Tab och bakåt med Skift + Kommando Ctrl +Tab.  
Redigera - AutoText  
Ordkomplettering  
Undantagslistan i AutoKorrigering  
Du kan återställa ett ord som korrigerats av AutoKorrigeringen med Ångra-funktionen.  
Ordet läggs då till i undantagslistan för AutoKorrigeringen, under förutsättning att funktionen "Lägg till automatiskt" är aktiverad i dialogrutan AutoKorrigering. (Förinställningen är att den är aktiverad.)  
Exempel  
AutoKorrigeringen korrigerar automatiskt ord som börjar med två stora bokstäver enligt standardinställningen.  
Men det kan vara meningen att produktnamn eller liknande ska skrivas så:  
Men AutoKorrigeringen gör automatiskt om det till "Est".  
Tryck på Kommando Ctrl +Z.  
Den automatiska ersättningen återställs och "ESt" läggs automatiskt till i undantagslistan i dialogrutan AutoKorrigering.  
Automatisk punktuppställning / numrering  
Om du aktiverar menyalternativet Format - AutoFormat - Under inmatningen känner %PRODUCTNAME automatiskt igen punktuppställningar och numreringar medan du skriver.  
Även romerska punktuppställningar resp. numreringar känns igen och fullföljs.  
Din numrering / punktuppställning kan börja på valfritt ställe i serien, den behöver med andra ord inte börja med t.ex. 1. eller I.  
Ett exempel på numrering med romerska siffror:  
Skriv ett I. (med punkt), följt av ett blanksteg och lite text.  
I stället för punkten kan du även välja en parentes.  
Tryck på returtangenten för att skapa ett nytt stycke.  
Det nya stycket börjar med II., romersk tvåa.  
Skriv lite text och tryck på returtangenten, så inleds nästa stycke med III. och så vidare.  
Du kan låta din romerska numrering börja med vilket tal som helst, t.ex. ci (motsvarar 101), följt av cii (102) och så vidare.  
Format - Numrering / Punktuppställning  
Stänga av automatiska ändringar  
I förinställningen korrigerar %PRODUCTNAME Writer ett stort antal vanliga skrivfel.  
Du kan ångra varje automatisk ändring direkt, t.ex. med Kommando Ctrl +Z.  
Här följer ställena i %PRODUCTNAME där du stänger av automatiska ändringar (och sätter på dem igen):  
Citatationstecken ersätts med typografiska anföringstecken  
Öppna ett textdokument.  
Välj Verktyg - AutoKorrigering / AutoFormat.  
Klicka på fliken Typografiska anföringstecken.  
Avmarkera Ersätt.  
Mening börjar alltid med stora bokstäver  
Öppna ett textdokument.  
Välj Verktyg - AutoKorrigering / AutoFormat.  
Klicka på fliken Alternativ.  
Avmarkera Börja varje mening med stor bokstav.  
Ord ersätts med ett annat ord  
Öppna ett textdokument.  
Välj Verktyg - AutoKorrigering / AutoFormat.  
Klicka på fliken Ersättning.  
Leta upp ordparet och radera det.  
Av tre lika tecken blir en hel linje  
Om du matar in tre av de följande tecknen i början av ett nytt stycke och sedan trycker på returtangenten blir det en hel linje av dem med olika styrka: - _ = * ~ #  
Öppna ett textdokument.  
Välj Verktyg - AutoKorrigering / AutoFormat.  
Klicka på fliken Alternativ.  
Avmarkera Använd inramning om du inte vill ha den här automatiska omvandlingen.  
Linjen är en inramning av det föregående stycket.  
Under Format - Stycke kan du redigera eller radera den.  
Automatisk rättstavningskontroll  
Alla ord som identifieras som felaktiga av rättstavningskontrollen stryks då under med en röd linje.  
Du kan klicka och samtidigt hålla ner Ctrl-tangenten med höger musknapp på de understrukna orden.  
Då visas en snabbmeny.  
På snabbmenyn finns det i många fall förslag på ord och du kan klicka på ett dem.  
Då ersätter förslaget ordet som är understruket med rött.  
Om du ersätter det felskrivna ordet via AutoKorrigering på snabbmenyn läggs ordparet in i AutoKorrigeringens ersättningstabell.  
Du kan öppna ersättningstabellen via Verktyg - AutoKorrigering / AutoFormat och fliken Ersättning.  
Om det understrukna ordet är rätt kan du lägga till det i en användarordlista med kommandot Lägg till.  
Utesluta ord från rättstavningskontrollen  
Markera orden.  
Öppna snabbmenyn till ett av orden.  
Välj Tecken.  
I dialogrutan Tecken klickar du på fliken Teckensnitt.  
Välj [inget] språk.  
Skapa användarordlistor  
Använda textblock som AutoText  
%PRODUCTNAME Writer innehåller en AutoText-funktion som gör att du kan sammanställa hela texter för brev, fax och valfria andra dokument genom att mata in förinställda förkortningar eller förkortningar som du själv definierar.  
Det finns följande möjligheter att infoga AutoText:  
Ange förkortningen för ett AutoText-block och tryck på F3.  
I programmet ingår flera färdiga AutoTexter:  
Om du t.ex. skriver BT och trycker på F3, infogas en typisk blindtext, ett stycke nonsenstext som kan hjälpa dig att bedöma utseendet på en sida som ska vara fylld med text (och andra objekt).  
Om du t.ex. skriver FN och trycker på F3, infogas en %PRODUCTNAME Math-formel med fortlöpande numrering i marginalen.  
Välj Redigera - AutoText.  
I dialogrutan AutoText finns det ett antal AutoTexter.  
Du kommer att märka att textblocken till och med kan innehålla grafik och tabeller.  
Klicka länge på ikonen AutoText på verktygslisten och välj en AutoText.  
Använd tipshjälpen med AutoComplete om du vill.  
Det finns anvisningar i %PRODUCTNAME -hjälpen.  
För muspekaren till textblocket som du vill infoga vid markörens position i texten.  
När du släpper musknappen infogas texten.  
Definiera AutoText  
Den kan innehålla formateringar och inbäddad grafik.  
Nu klickar du kort på ikonen Redigera AutoText på verktygslisten.  
Välj kategori (t.ex. "standard") i den stora listrutan, namnge det nya textblocket i textfältet och korrigera eventuellt förkortningen.  
Nu kan du spara textblocket med AutoText - Nytt och sedan stänga dialogrutan.  
AutoText i nätverk  
Du kan använda AutoTexter från olika kataloger.  
Ett exempel med en typisk nätverksinstallation av %PRODUCTNAME:  
I en katalog på servern kan företagets skrivskyddade AutoTexter stå medan du skriver och läser dina egna, användardefinierade AutoTexter i ditt eget filområde.  
Välj Verktyg - Alternativ - %PRODUCTNAME - Sökvägar.  
Dubbelklicka på posten AutoText.  
Här är redan två sökvägar angivna.  
Den första sökvägen gäller AutoTexterna från serverinstallationen, den andra sökvägen AutoTexterna från din userkatalog.  
Om två AutoTexter från olika kataloger har samma namn använder %PRODUCTNAME AutoTexten från din userkatalog.  
Skriva ut AutoTexter  
Då listas alla namn och förkortningar för AutoTexterna i ett nytt textdokument.  
Välj Verktyg - Makro..., dubbelklicka på "Gimmicks" i listan till höger i dialogrutan Makro, markera "AutoText "och klicka på Kör.  
Redigera - AutoText  
Ordkomplettering  
Räkna med formler som står i text  
Om det redan finns en matematisk formel i texten kan du kopiera beräkningen av resultatet till texten utan att använda formellisten:  
Markera den matematiska formeln i texten som inte får innehålla någonting annat än siffror, räknekommandon och eventuella valutabeteckningar.  
Exempel:  
12 + 24 * 2  
Tryck på Kommando Ctrl + (plustecknet), eller välj Verktyg - Beräkna.  
Resultatet av beräkningen finns nu i urklippet.  
Tryck på Kommando Ctrl +V, eller välj Redigera - Klistra in.  
I exemplet infogas 60.  
Om formeln fortfarande är markerad när resultatet klistras in ersätter det formeln.  
Beräkna summor av tabellceller  
Foga in en tabell med flera rader i ett tomt textdokument (Infoga - Tabell).  
Lämna den nedersta cellen i kolumnen tom.  
Klicka sedan på ikonen Summa på tabellobjektlisten.  
På inmatningsraden står summaformeln med cellerna som står ovanför den här cellen, i form av en lista med summander.  
Mellan de enskilda summanderna finns listavgränsaren i form av ett lodstreck (_BAR_).  
Bekräfta genom att trycka på returtangenten eller klicka på Överta på formellisten.  
Summan visas i den nedersta cellen.  
När du ändrar talen i texttabellen uppdateras summan automatiskt.  
Om du t.ex. vill formatera talen i valutaformat, markerar du motsvarande celler och väljer Talformat på snabbmenyn.  
Dialogrutan Talformat visas, där du kan välja alla format.  
Räkna med tabeller i textdokument  
Du kan göra beräkningar i tabeller i %PRODUCTNAME Writer.  
Vid beräkningar som går utanför den aktuella tabellen fungerar tabellnamnet som entydig identifikation av tabellen.  
Om du t.ex. multiplicerar den första cellen i Tabell1 med den första cellen i Tabell2 och vill spara resultatet i cell A2 i den aktuella tabellen, placerar du markören i cell A2 i den aktuella tabellen, trycker på F2 och skriver sedan följande kommando på beräkningsraden:  
=<Tabell1.A1> * <Tabell2.A1>  
Med hjälp av Navigationslisten kan du förflytta dig mellan tabellformlerna i dokumentet.  
Om det finns en referens till en ogiltig tabellcell i en tabellformel, visas meddelandet "**Felaktigt uttryck**" i cellen.  
Ogiltiga tabellceller är raderade celler eller celler som innehåller fel.  
Om du vill addera innehållet i cellerna B1:B10 i Tabell1 och få resultatet i den encelliga Tabell2, som ska placeras någonstans i texten, gör du så här:  
Skapa texten och Tabell1.  
Skriv den text där resultatet ska visas.  
Infoga nu en ram (med menykommandot Infoga - Ram).  
I dialogrutan Ram väljer du förankringen Vid tecken och tar bort inramningen.  
Avmarkera ramen genom att klicka utanför den, och klicka sedan mitt i den som när du ska skriva text i den.  
Ramen får inte vara markerad; däremot ska textmarkören stå inuti ramen.  
Infoga den encelliga Tabell2 i ramen (Infoga - Tabell).  
Välj en rad och en kolumn och klicka på OK.  
Inmatningsmarkören står i Tabell2.  
Definiera nu en beräkningsformel genom att skriva ett likhetstecken.  
Formellisten visas.  
Markera de celler där posterna, som ska summeras i formeln, står i Tabell1 genom att hålla ner musknappen och föra muspekaren från den första till den sista cellen.  
Formeln för beräkning av summan av cellerna B1 till B10 lyder: =<Tabell1.B1:B10>  
Stäng formeln genom att klicka på ikonen Överta på formellisten.  
Resultatet visas i Tabell2.  
Om du ändrar de summerade talen kan du uppdatera resultatet genom att trycka på funktionstangenten F9.  
I stället för att först infoga ramen och sedan infoga en tabell i den, kan du först infoga en encellig tabell, markera den - i det här fallet går det bara med tangentkombinationen Kommando Ctrl +A - och sedan klicka på ikonen Infoga - Ram.  
Ramen omger då automatiskt tabellen (detta fungerar för övrigt även för textavsnitt).  
Nu kan du ställa in förankringen Vid tecken, klippa ut det hela till urklippet och klistra in det på önskad plats, ta bort inramningarna från ram och tabell och göra fler inställningar.  
Beräkning i text  
Placera markören på det ställe i texten där resultatet skall fogas in.  
Visa formellisten genom att trycka på F2.  
Mata in den önskade formeln, t.ex. (4+6 )*100.  
Infoga resultatet genom att trycka på returtangenten eller klicka på ikonen Överta.  
Om du ska genomföra en mer komplicerad beräkning kan du använda ikonen Formel.  
När du klickar på den öppnas en undermeny där du väljer en formel.  
Formeln infogas vid markörens position på formellisten.  
Du kan växla mellan att ange formler och värden med tangentbordet eller med ikonen Formel.  
Som ett exempel på en litet mer komplicerad beräkning i texten beräknar vi medelvärdet av tre tal.  
Öppna formellisten med F2.  
Öppna undermenyn till ikonen Formel.  
Välj Medelvärde under Statistiska funktioner.  
På inmatningsraden står det nu =mean.  
Mata in det första talet, och sedan listavgränsaren (_BAR_), d.v.s. ett lodrätt streck.  
Mata in det andra talet, ytterligare en listavgränsare och sedan det tredje talet.  
På inmatningsraden kan det nu t.ex. stå: =mean 12_BAR_ 22 _BAR_34  
Tryck på returtangenten så visas resultatet i texten.  
Det har infogats i form av ett fältkommando.  
Om du vill redigera ett fältkommando dubbelklickar du på det.  
Beräkningar i flera tabeller  
Foga in två tabeller med flera rader och kolumner i ett textdokument.  
Men låt minst en cell vara tom.  
Tabellerna kallas automatiskt för "Tabell1" och "Tabell2 ".  
Du kan också ge en tabell ett eget namn (Format - Tabell, fliken Tabell, textfältet Namn).  
Använd inga andra tecken än bokstäver och siffror i namnet.  
Placera markören i en tom cell.  
Tryck på F2.  
Formellisten visas.  
Skriv SUM som exempel.  
Nu kan du klicka i cellerna med tal i båda tabellerna.  
Sedan klickar du på nästa cell med ett tal.  
Slutligen klickar du på ikonen Överta på formellisten.  
Om du t.ex. vill summera de båda första cellerna i varje tabell och summan skapas i Tabell2, är formeln =sum <Tabell1.A1> + <A1>.  
Räkna i ett textdokument  
Du kan göra beräkningar i textdokument, både i löpande text och i tabeller som du har skapat i textdokumenten.  
Formellisten visas om du trycker på funktionstangenten F2 i en tabellcell eller någonstans i texten.  
I en tabell räcker det om du skriver ett likhetstecken.  
Detta signalerar att du vill mata in en matematisk formel.  
Du döljer formellisten igen genom att trycka på F2 eller på Esc.  
Så här räknar du direkt i texten  
Du skriver t.ex. följande text: "$10000 per år, det är $i månaden."  
Placera markören på den plats där du vill infoga resultatet och tryck på F2.  
Formellisten visas och markören är redan placerad där.  
Mata in 10000 / 12 och tryck på Retur.  
Resultatet av beräkningen infogas i texten.  
Numrera bildtexter efter kapitel  
Om du vill numrera alla illustrationer i dokumentet kapitelvis så att illustrationerna i det första kapitlet t.ex. har bildtexterna "Illustration 1.1", "Illustration 1.2" o.s.v., och bilderna i det andra kapitlet "Illustration 2.1", "Illustration 2.2 "o.s.v., gör du så här:  
Dela upp dokumentet i kapitel, om du inte redan har gjort det.  
Välj Verktyg - Kapitelnumrering... och tilldela kapitelöverskrifterna, som du t.ex. har formaterat med styckeformatmallen "Överskrift 1", en numrering.  
I listrutan väljer du mallen "Överskrift 1" som styckeformatmall, och i listrutan nedanför väljer du alternativet "1, 2, 3 "under Nummer.  
Välj den första illustrationen som du vill numrera.  
Välj Infoga - Bildtext...  
I den dialogruta som nu visas väljer du posten Illustration som kategori och "Arabiska siffror (1 2 3)" som numrering.  
Här kan du också skriva bildtexten.  
Klicka på Alternativ.  
I dialogrutan Sekvensalternativ kan du bestämma hur den kapitelvisa numreringen ska göras.  
I exemplet väljer du alternativ "1" under Nivå och anger ett skiljetecken för den kapitelvisa numreringen.  
Bekräfta med OK.  
Om du nu slutligen bekräftar dialogrutan Bildtext med OK numreras illustrationen efter sitt kapitel.  
Gör likadant med alla andra illustrationer i dokumentet.  
Alla illustrationer på en och samma kapitelnivå numreras löpande.  
I dialogrutan Sekvensalternativ anger du mellan vilka kapitelnivåer numreringen ska växla.  
Under Verktyg - Alternativ - Textdokument - Allmänt kan du markera rutan Bildtext - Automatiskt.  
Om du nu klickar på kommandoknappen bredvid Objekturval visas dialogrutan Bildtext.  
Här kan du definiera att t.ex. alla illustrationer ska få en automatisk bildtext i textdokument i framtiden.  
Bildtexter och nummersekvenser  
I textdokument kan du skapa separata bildtexter med löpande numrering för illustrationer, tabeller och ritobjekt.  
Du kan definiera ett valfritt antal egna nummersekvenser.  
Bildtexterna är kopplade till illustrationerna, tabellerna eller ritobjekten i en ram.  
Markera ramen om du flyttar objektet.  
Definiera bildtexter  
Markera illustrationen eller objektet eller placera markören i den tabell för vilken du vill infoga en bildtext.  
Välj Infoga - Bildtext.  
Dialogrutan Bildtext visas.  
I dialogrutan ser du i en förhandsvisning hur bildtexten ser ut.  
Du kan lägga till fler texter i fältet Bildtext.  
Klicka på OK.  
Om du vill ha ett tabbsteg mellan den automatiska bildtexten av typen "Illustration 1" och din tilläggstext, kan du infoga detta i dokumentet i efterhand.  
Tryck på Ctrl+Tabb för att infoga en tabb i början av ett stycke.  
Styckeformatet för den automatiskt infogade bildtexten hämtas från styckeformatmallen "Illustration", "Tabell", "Teckning" eller "Text ".  
De här styckeformatmallarna baserar alla på styckeformatmallen "Bildtext".  
Om du alltså vill att alla bildtexter alltid ska visas i grönt, behöver du bara göra motsvarande ändring i styckeformatmallen "Bildtext" i Stylist.  
Använd vyalternativet "Alla mallar" eller hierarkisk visning i Stylist.  
Redigera eller radera bildtext  
Bildtexten är normal text som står tillsammans med objektet i en gemensam ram.  
Redigera bildtexten som normal text.  
Radera bildtexten som normal text.  
Infoga objekt i en nummersekvens  
Utöka den automatiska nummersekvensen "Illustration" på följande sätt:  
Tilldela stycket styckeformatmallen "Illustration".  
Styckets innehåll kan bestå av ordet "Illustration" med ett följande blanksteg.  
Öppna sedan dialogrutan Fältkommandon, t.ex. med Kommando Ctrl +F2.  
Välj fälttypen "Nummersekvens" under fliken Variabler.  
Under Urval väljer du "Illustration".  
Klicka på Infoga och stäng dialogrutan.  
Om du vill flytta illustrationer med deras bildtexter för hand så att ordningsföljden ändras, måste du eventuellt uppdatera visningen av nummer med F9.  
Sidformatmall från markering  
Ofta behövs en ny sidformatmall, t.ex. därför att sidhuvudet ska ändras vid kapitelväxling.  
Sidhuvudet är kopplad till sidformatmallen.  
Eftersom attributen i formatmallen ofta inte ändras för övrigt, bör en sådan formatmall skapas via funktionen "Ny mall från markering" i Stylist.  
Den nya mallen övertar då automatiskt alla mallens attribut från sidan där markören står.  
Du har skapat en sidformall med en viss text i sidhuvudet och skrivit flera sidor.  
På de följande sidorna ska en annan text finnas i sidhuvudet.  
Växla till Sidformatmallar i Stylist.  
Den nya sidformatmallen tilldelar du de följande sidorna.  
Välj kommandot Infoga - Manuell brytning.  
Välj alternativet Sidbrytning i området Typ och välj den nya mallen i listrutan.  
Skriv den nya texten i sidhuvudet på en av de nya sidorna.  
Den gäller då för alla sidor med den här sidformatmallen.  
Kapitelnumrering  
På meny Verktyg - Kapitelnumrering kan du låta numrera dina överskrifter automatiskt.  
I förinställningen är den översta nivån i kapitelnumreringen tilldelad styckeformatet "Överskrift 1".  
Om du väljer en numreringstyp i kombinationsfältet Nummer, sätts ett löpande nummer framför alla stycken som har formatet "Överskrift 1" i ditt dokument.  
Om du har gjort egna styckeformatmallar som du vill använda för överskrifter, kan du tilldela de enskilda nivåerna mallarna i den här dialogrutan.  
Om du t.ex. har gjort en styckeformatmall som heter "Head1" och som används för överskrifterna på nivå 1, väljer du 1 under Nivå och Head1 i kombinationsfältet Styckeformatmall.  
Klicka på OK.  
Nu listas alla stycken som formateras med Head1 i Navigator under "Överskrifter".  
Du kan placera om kapitlen i Navigator om du vill ändra deras ordning eller nivå i hierarkin och på så sätt även numreringen:  
Klicka på en av ikonerna Kapitel uppåt, Kapitel nedåt, En nivå upp och En nivå ner, eller  
flytta kapitelöverskriften i Navigator med musen.  
Numreringen av alla berörda kapitel anpassas automatiskt.  
Villkorlig text för sidantal  
Hur får man ordet "Sida" att skrivas korrekt i visningen av sidantal i ett textdokument (alltså "Sida "eller "Sidor")?  
För att göra skrivsättet av ordet "Sida" oberoende av det faktiska sidantalet finns fältkommandot Villkorlig text.  
Gör på följande sätt:  
1.  
Placera markören på det ställe i dokumentet där sidor sidnumret skall anges.  
2.  
Välj meny Infoga - Fältkommando - Sidantal.  
Sidantalet infogas i dokumentet.  
Foga in ett blanksteg direkt efter.  
3.  
Välja meny Infoga - Fältkommando - Andra.  
Välj fliken Funktioner och klicka sedan på Villkorlig text under Fälttyp.  
4.  
I fältet Villkor matar du in: "Page > 1" (utan citationstecken).  
I fältet Så matar du in: "Sidor" I fältet Annars matar du in: "Sida "  
5.  
Klicka på Infoga för att infoga fältkommandot i dokumentet och sedan på Stäng för att avsluta fältkommandodialogen.  
Beroende på antalet sidor används nu det korrekta skrivsättet.  
Uppdatering av visningen sker med tangenten (F9).  
Villkorlig text  
Anta att du t.ex. vill att ett visst stycke bara ska visas i dokumentet om ett särskilt villkor är uppfyllt, och i annat fall att ett annat stycke ska visas.  
Ett bra exempel är ett påminnelsebrev, som vid tredje påminnelsen innehåller andra formuleringar än vid den första.  
Detta kan du uppnå med fältkommandot "Villkorlig text".  
Högre upp i ditt påminnelsebrev finns det en rad "1:a påminnelsen" till "3:e påminnelsen ".  
Talet anger du som användardefinierad variabel i ett fältkommando.  
Placera markören på det ställe där det löpande numret 1 till 3 ska visas i dokumentet.  
Öppna dialogrutan Fältkommando (t.ex. med Kommando Ctrl +F2) och växla till fliken Variabler.  
Välj fälttypen "Sätt variabel".  
Ange ett namn för den nya variabeln i textfältet Namn, t.ex. "Påminnelse".  
Välj Text som variabelformat.  
Ange värdet 1 i textfältet Värde och klicka på Infoga.  
Placera nu markören på det ställe i texten där den villkorliga texten ska infogas.  
Dialogrutan Fältkommando finns kvar på bildskärmen tills du stänger den.  
Välj fälttypen "Villkorlig text" under fliken Funktioner.  
Nu ska du ange ett villkor.  
I vårt fall lyder det Påminnelse EQ "3".  
De operatorer som får användas i den här typen av logiska sökningar hittar du i en lista över operatorer i %PRODUCTNAME -hjälpen.  
Talet 3 står här inom citattecken, vilket innebär att du inte söker efter det numeriska värdet utan efter texttecknet.  
När variablerna definierades var ju posten Text markerad - om du hade markerat Tal där, skulle du kanske nu bli förvånad över de decimaler som visas i standardformatet för tal. "1,00 påminnelse" som överskrift ser något ovanligt ut.  
I stället för format Text kan du välja formatet "1234567", för att bara visa heltal.  
Under Så skriver du den text som ska infogas om det är den tredje påminnelsen.  
Under Annars skriver du den text som ska visas i de andra fallen.  
Det finns ingen begränsning för textens längd.  
Om du vill kan du kopiera texten direkt från ett dokument till textinmatningsfältet.  
Klicka på Infoga och stäng dialogrutan.  
Vid behov kan du visa eller dölja fältkommandona genom att trycka på Kommando Ctrl +F9.  
Om du i stället för en "1:a påminnelse" vill skriva en "2:a "eller "3:e påminnelse", så placerar du textmarkören direkt framför fältkommandot med innehållet "1" och väljer kommandot Redigera - Fältkommando, eller så dubbelklickar du på det gråmarkerade fältkommandot.  
Ange sedan tecknet "2" eller "3 "i stället för "1" i dialogrutan och stäng den sedan.  
Du ser texten till den sista påminnelsen i dokumentet.  
Denna tangent uppdaterar alla beräkningar i ett dokument.  
Ta bort ord från användarordlista  
Välj Verktyg - Alternativ - Språkinställningar och sedan Lingvistik.  
Markera användarordlistan och klicka på Redigera.  
Nu visas dialogrutan Redigera användarordlista där du kan söka igenom en lista i alfabetisk ordning.  
Markera ordet och klicka på Radera.  
Flytta textavsnitt i dokument  
Markera texten som du vill flytta.  
Peka på den markerade texten, tryck sedan på musknappen och håll ner den.  
Dra bort musen en bit.  
Du ser en symbol bredvid pekaren som visar att det markerade området flyttas.  
Markören följer pekaren och antyder målet för förflyttningen.  
Muspekare - form  
Betydelse  
Flytta  
Kopiera  
Om du inte vill flytta texten utan bara kopiera den, håller du ner Kommando Ctrl -tangenten medan du gör dra-och-släpp.  
Muspekaren visar detta med ett plustecken.  
Du kan trycka ner och släppa Kommando Ctrl -tangenten så ofta du vill - det är tillståndet som råder när man släpper musknappen som gäller.  
Byta sidformatmall på jämna och ojämna sidor  
Om du t.ex. vill ha annat innehåll i sidhuvudena och sidfötterna på jämna sidor (vänstersidor) än på ojämna sidor (högersidor) definierar du det i sidformatmallarna.  
Använd olika siformatmallar för vänster - och högersidor.  
Definiera att en högersida kommer som nästa formatmall efter en vänstersida och att en vänstersida kommer efter en högersida.  
Öppna Stylist.  
Klicka på ikonen Sidformatmallar i Stylist.  
Klicka på sidformatmallen Vänstersida och öppna sedan snabbmenyn.  
Välj kommandot Ändra.  
Dialogrutan Sidformatmall: Vänstersida  
Klicka på fliken Administrera.  
I fältet Nästa formatmall väljer du Högersida.  
På samma sätt ändrar du mallen Högersida så att den har Vänstersida som nästa formatmall.  
Tilldela den första sidan i dokumentet sidformatmallen Högersida.  
Det gör du t.ex. genom att sätta markören på den första sidan i dokumentet och sedan dubbelklicka på sidformatmallen Högersida i Stylist.  
På statuslisten visas alltid vilken sidformatmall som gäller.  
Om du vill ha en titelsida som inte innehåller något sidhuvud eller någon sidfot, gör du så här:  
Ändra sidformatmallen Första sidan så att den har Vänstersida som nästa formatmall.  
Tilldela din titelsida sidformatmallen Första sidan.  
Dialogrutan Infoga brytning  
Omvandla fältkommando till text  
Du vill omvandla det här fältkommandot till normal text.  
Placera markören bredvid fältkommandot.  
Skriv av innehållet i fältkommandot (i det här exemplet datumet).  
Radera fältkommandot.  
Alternativt använder du urklippet på följande sätt:  
Markera fältkommandot (i det här exemplet datumet).  
Klipp ut fältkommandot till urklippet, t.ex. med Redigera - Klipp ut.  
Klicka länge på ikonen Klistra in på funktionslisten.  
I undermenyn väljer du Oformaterad text.  
Textinnehållet i fältkommandot klistras in.  
Redigera - Klistra in innehåll  
Infoga datum fast eller variabelt.  
Så här infogar du ett variabelt datum i %PRODUCTNAME Writer.  
Öppna meny Infoga - Fältkommando - Andra... och välj fältkommandot Datum under fliken Dokument.  
Fältkommandot för ett variabelt datum kommer att visa aktuellt datum enligt systemtiden varje gång dokumentet öppnas och när fältkommandona uppdateras.  
I motsats till detta infogar fältkommandot Datum (fast) ett datum som alltid motsvarar det datum som gällde när det infogades.  
När dokumentet öppnas eller uppdateras en annan dag förblir det fasta datumet oförändrat.  
Skapa inmatningsfält i text  
Så skapas ett textdokument med inmatningsfält där markören hoppar direkt till nästa fält.  
I %PRODUCTNAME Writer finns fältkommandot Inmatningsfält (på meny - Infoga - Fältkommando - Andra - flik Funktioner).  
De här inmatningsfälten kan du placera på de ställen i dokumentet där användaren skall infoga variabel text.  
Via tangentkombinationen Ctrl+Skift+F9 eller genom att dubbelklicka på fältkommandot kan du öppna en dialogruta där du kan ändra innehållet.  
Söka användardata i villkor  
I fältformler eller villkor har du även åtkomst till användardata.  
Användardata är strängar som du kan jämföra med följande operatorer:  
Operator  
Betydelse  
== eller EQ  
är lika med  
!= eller NEQ  
är inte lika med  
Det finns fler operatorer i %PRODUCTNAME -hjälpen.  
Så här döljer du ett området för en användare  
Markera texten som användaren "Andersson" inte ska se.  
Välj kommandot Infoga - Område.  
Markera fälten Dölj och Med villkor.  
Skriv in villkoret i textfältet:  
user_lastname == "Andersson"  
Klicka på Infoga och spara dokumentet.  
Om den nämnda användaren öppnar textdokumentet, kan han eller hon inte se området.  
I Navigator visas namnet på området.  
Om en annan användare öppnar samma textdokument, kan han / hon se området.  
Följande tabell innehåller användarvariablerna.  
Användarvariabel  
Betydelse  
user_firstname  
Förnamn  
user_lastname  
Efternamn  
user_initials  
Initialer  
user_company  
Företag  
user_street  
Gatuadress  
user_country  
Land  
user_zipcode  
Postnummer  
user_city  
Ort  
user_title  
Titel  
user_position  
Befattning  
user_tel_work  
Telefon - arbetet  
user_tel_home  
Telefon - privat  
user_fax  
Faxnummer  
user_email  
E-postadress  
user_state  
Delstat  
Använda fältkommandon  
Via fältkommandon kan du t.ex. infoga aktuellt datum, aktuellt sidnummer, dokumentets totala antal sidor, korshänvisningar till andra ställen i texten, innehållet i vissa databasfält från en databas och ett stort antal andra variabler, d.v.s. värden som ändras, i dokumentet.  
Den största fördelen med fältkommandon ligger i att %PRODUCTNAME övervakar fältinnehållets utseende och eventuellt anpassar det till dokumentets aktuella redigeringsstatus.  
Hur visas fältkommandon?  
Fältkommandon består i princip av elementen Fältnamn och Fältinnehåll.  
Med menykommandot Visa - Fältkommandon kan du växla mellan visning av fältnamn och fältinnehåll.  
Om du har markerat rutan Fixera innehåll, förses fältnamnet i fråga med tillägget "fix".  
Fältkommandonas bakgrund i färg kan du sätta på och stänga av under Verktyg - Alternativ - Textdokument - Vy med funktionen Bakgrund Fält.  
Du kan även sätta på och stänga av bakgrunden med menykommandot Visa - Markeringar.  
Vid HTML-import och -export gäller särskilda %PRODUCTNAME -definierade taggar för fältkommandon.  
Vilka egenskaper har fältkommandon i dokumentet?  
Det finns olika typer av fältkommandon, som uppträder på olika sätt, beroende på vilken funktion de har:  
De flesta fälten används för att lägga till variabelt innehåll och infoga det i aktuell form i dokumentet.  
Det kan vara dokumentinformation eller databasinnehåll.  
Några fält utför en åtgärd när man klickar på dem med musen.  
Dessa fält känner man igen på att de antar formen av en hand, när man för pekaren över dem.  
Åtgärderna kan vara olika definierade beroende på fälttyp.  
Du har följande alternativ:  
Fälttyp  
Egenskap  
Platshållare  
Genom att klicka öppnar du en dialogruta där du kan infoga det objekt för vilket platshållaren har satts.  
Infoga referens  
Du placerar markören på den satta referensen genom att klicka.  
Utför makro  
Du startar makrot genom att klicka.  
Inmatningsfält  
Genom att klicka öppnar du en dialogruta där du kan redigera innehållet.  
Vid några fälttyper visas en kort hänvisningstext, namnet eller fältets värde, om du placerar markören på detta fält.  
Du anger de visade hänvisningarna, beteckningarna eller värdena i motsvarande textfält i dialogrutan Fältkommandon.  
Detta gäller för variabler, databasfält, användardefinierade fält och fält av typen Platshållare, Dold text samt "Infoga referens".  
Hur uppdateras fältkommandon?  
Om du vill uppdatera fältinnehållen räcker det i de flesta fall att du trycker på funktionstangenten F9.  
Vid infogade databasfält markerar du fältkommandot och trycker sedan på F9.  
Om du vill uppdatera alla fältkommandona i dokumentet, väljer du menykommandot Redigera - Markera allt eller Kommando Ctrl +A och trycker sedan på F9.  
Redigera text med FontWork  
Du kan skapa grafiska texteffekter med programmodulen FontWork.  
Gör så här:  
1.  
Öppna utrullningslisten Ritfunktioner på verktygslisten och klicka på ikonen Text.  
2.  
Rita upp en textram och skriv sedan in en text, till exempel "FontWork".  
3.  
Välj Format - FontWork.  
Du ser FontWork-fönstret där du väljer effekter:  
4.  
Klicka på ikonen uppe till vänster med halvcirkeln som är böjd uppåt.  
Texten visas i bågform.  
5.  
Bland alternativen för skugga klickar du på Lodrätt.  
Ställ in värdet "2,00mm" i fältet med rotationsknapparna för att öka skuggan på X-axeln.  
Texten ser redan nu nästan ut som på bilden.  
6.  
Du behöver bara dubbelklicka på texten, redigera den och sedan klicka utanför objektet.  
7.  
Om du markerar FontWork-objektet genom att klicka med musen, ser du åtta handtag.  
Du kan dra en av dessa handtag med musen och därigenom ändra hela objektets storlek och form.  
Det färdiga objektet kan du kopiera via urklippet och klistra in i andra dokument, ändra storleken där och så vidare.  
Format - FontWork  
Infoga följande sidas sidnummer  
Infoga först en sidfot via Infoga - Sidfot.  
Placera sedan markören i sidfoten och välj Infoga - Fältkommando - Andra....  
Klicka på fliken Dokument och välj fälttypen "Sida" och under Urval "Nästa sida ".  
Välj "Som sidformatmallen" under Format och klicka sedan på Infoga för att infoga fältkommandot i sidfoten för det aktuella dokumentet.  
I ditt dokument kommer nu sidnumret på nästa sida att visas på varje sida, utom på den sista sidan naturligtvis.  
Om dessutom ordet "Sida" ska visas framför sidnumret infogar du helt enkelt ytterligare ett fältkommando av samma typ, men i ett annat format:  
Sätt markören framför fältkommandot som du precis har infogat och öppna dialogrutan Fältkommando igen.  
Välj ett fältkommando av typen "Sida" igen, välj "Nästa sida "igen under Urval och sedan "Text" under Format.  
I textfältet Värde kan du nu mata in en text som ska visas när det finns en sida till.  
Mata in "fortsätter på sida" (med ett mellanslag) och klicka sedan på Infoga.  
I stället för "sida" kan du givetvis även mata in andra tecken, t.ex. "... / "för att markera att numret på följande sida står här.  
Infoga sidnummer i sidfot  
Infoga en sidfot.  
Välj Infoga - Sidfot och välj på undermenyn för vilken sidformatmall du vill ha sidfoten.  
Markören står nu i sidfoten.  
Välj Infoga - Fältkommando - Sidnummer.  
Du ser sidnumret som fältkommando i sidfoten.  
Markera sidnumret och klicka på ikonen Centrerat på objektlisten.  
Om du vill ha sidfotstexten i form av "Sida 9 av 12", gör du så här:  
Skriv texten "Sida" före fältkommandot och "av" efter fältkommandot.  
Välj Infoga - Fältkommando - Sidantal.  
Infoga och redigera fotnoter  
Du kan infoga en fotnot på två sätt, med hjälp av en ikon eller med en dialog.  
Så här infogar du en fotnot med en ikon  
1.  
Placera markören på det ställe i texten där fotnotsankaret ska visas.  
2.  
Öppna utrullningslisten Infoga på verktygslisten.  
3.  
Klicka på ikonen Infoga fotnot direkt.  
Så här infogar du en fotnot med en dialogruta  
Placera markören på det ställe i texten där fotnotsankaret ska visas.  
Välj Infoga - Fotnot.  
Dialogrutan Infoga fotnot öppnas.  
När du infogar en fotnot med ikonen används en automatisk fotnotsnumrering, medan dialogrutan Infoga fotnot innehåller möjligheter att göra inställningar för fotnoten.  
Information om hur du arbetar med fotnoter  
Om du vill redigera texten i en fotnot, klickar du på den och ändrar den.  
Du kan hoppa från fotnotsområdet till fotnotsankaret i texten med Page Up-tangenten.  
Om du vill redigera egenskaperna för en infogad fotnot, placerar du markören omedelbart framför fotnotstecknet i dokumentet och väljer Redigera - Fotnot eller dubbelklickar omedelbart framför fotnotstecknet.  
I dialogrutan Fotnotsinställning som du öppnar via Verktyg - Fotnoter gör du allmängiltiga inställningar som ska användas automatiskt för fotnoter i dokumentet.  
Formateringen av fotnotsområdet görs via sidformatmallen.  
Välj Format - Sida... - Fotnot.  
På sidor med flera kolumner infogas fotnoten i kolumnen där fotnotsankaren finns.  
Du kan även hoppa från fotnotsankaret till fotnoten med musen.  
Muspekaren byter utseende när du pekar på fotnotsankaret.  
Avstånd mellan fotnoter  
Om du vill ha ett större avstånd mellan enskilda fotnoter eller slutnoter kan du lägga till en osynlig (vit) linje som undre inramning till motsvarande styckeformat:  
Placera markören i en fotnot.  
Öppna Stylist.  
Klicka på styckeformatmallen som ska ändras (Fotnot).  
Öppna snabbmenyn och välj Ändra.  
Ge båda färgen vitt.  
I området Avstånd till innehåll tar du bort markeringen i rutan Synkronisera.  
Höj värdet för det övre och undre avståndet.  
Klicka på OK.  
Format - Stycke - Inramning  
Använda samlingsdokument och deldokument  
Du kan välja mellan att skapa ett nytt tomt samlingsdokument (Arkiv - Nytt - Samlingsdokument) eller att skapa ett samlingsdokument utifrån ett befintligt dokument via Arkiv - Skicka - Skapa samlingsdokument.  
Du öppnar ett nytt samlingsdokument genom att välja Arkiv - Nytt - Samlingsdokument.  
Det nya samlingsdokumentet öppnas som ett tomt textdokument och samtidigt visas Navigator i samlingsläge.  
Navigator i samlingsläge har bland annat funktioner som du använder för att navigera och redigera.  
Du laddar ett dokument för redigering genom att dubbelklicka på det i Navigator.  
Lägg märke till filnamnstillägget ".sgl" när du öppnar ett befintligt samlingsdokument. "Normala "%PRODUCTNAME Writer-dokument har filnamnstillägget ".sxg".  
Ett exempel på ett samlingsdokument finns bland %PRODUCTNAME -exemplen.  
Lägg in text, t.ex. för överskrifter, eller infoga deldokument genom att klicka på ikonen Infoga och välja önskad post Text eller Fil.  
I så fall anger du först ett namn och var det ska sparas.  
Styckeformatmallar som du definierar och använder i deldokumenten tas automatiskt upp i samlingsdokumentet.  
Om du sparar samlingsdokumentet efter det är de här formatmallarna tillgängliga i alla delar av samlingsdokumentet.  
Formatmallar som har definierats i samlingsdokumentet har högre prioritet än formatmallarna med samma namn i deldokumenten.  
Det bästa är att basera alla deldokument och själva samlingsdokumentet på en och samma dokumentmall.  
Om du behöver en ny formatmall i dokumenten infogar du den bara i dokumentmallen och laddar samlingsdokumentet på nytt.  
Du kan automatiskt överföra den nya formatmallen till alla dokument.  
Om alla deldokument ska börja på en ny sida (kanske t.o.m. alltid på en ny högersida) kan du arbeta med sidformatmallar.  
Det finns en färdig sidformatmall som heter "Höger sida" som du t.ex. kan koppla till styckeformatmallen "Överskrift 1 ".  
Om du tilldelar styckeformatmallen "Överskrift 1" en sidbrytning hamnar alla "Överskrift 1 "alltid överst på en högersida.  
Som nästa formatmall tilldelar du sidformatmallen "Högersida" "Vänstersida "och tvärtom.  
När markören står i en text i ett samlingsdokument är posten Text nedtonad eftersom texter som står i följd alltid sammanfogas till en enda text.  
Du kan infoga ny text mellan enskilda infogade dokument.  
Men du kan lätt ändra ordningsföljden genom att dra och släppa eller genom att klicka på ikonerna Flytta nedåt respektive Flytta uppåt.  
Dokument infogas som skyddade områden i samlingsdokumentet.  
Men du kan bläddra i dokumenten för att läsa dem.  
Förteckningarna omfattar automatiskt alla deldokument.  
Om du ändrar ett eller flera deldokument när du har skapat en förteckning måste du uppdatera förteckningarna i samlingsdokumentet.  
Klicka på ikonen Uppdatera i Navigator för samlingsdokument och välj vad du vill uppdatera på undermenyn.  
Referenser fungerar mellan samlingsdokument och deldokument samt inom deldokument om de är enhetliga i alla dokument som finns med.  
Om bilderna i ett deldokument är numrerade från "Bild 1" till "Bild 10 "ska bilderna fortsätta med "Bild 11" i nästa deldokument.  
Om du vill kan du spara samlingsdokumentet med alla delar som ett %PRODUCTNAME Writer-dokument.  
Välj Arkiv - Spara som och välj ett "normalt" %PRODUCTNAME Writer-format i listrutan Filtyp.  
När du skriver ut ett samlingsdokument skrivs alla deldokument, texter och förteckningar ut.  
Håll muspekaren över den aktuella posten i Navigator.  
Sökvägen till originaldokumentet visas i ett litet fönster.  
Om filen inte finns kvar på den ursprungliga platsen visas, förutom sökvägen, meddelandet Filen har ej hittats i rött.  
Information om sidhuvuden och sidfötter  
Sidhuvuden och sidfötter är alltid kopplade till sidformatmallen.  
Samtliga sidor med samma sidformatmall har automatiskt samma sidhuvuden och sidfötter.  
Du kan infoga variabla innehåll i textdokument, t.ex. sidnummer och kapitelöverskrifter, med hjälp av fältkommandon i sidhuvuden och sidfötter.  
Om du vill ha ytterligare skillnader i sidhuvudenas och sidfötternas innehåll är det bäst att skapa olika sidformatmallar och tilldela sidorna dem.  
Under Infoga - Sidhuvud eller Infoga - Sidfot kan du välja för vilken sidformatmall du vill infoga eller ta bort sidhuvuden eller sidfötter.  
I dialogrutan Format - Sida kan du också välja om du vill ha sidhuvuden eller sidfötter i den aktuella sidformatmallen.  
Här finns det också en ruta som heter Samma innehåll till höger / vänster och om den inte är markerad, kan du formatera olika sidhuvuden och sidfötter på vänster - och högersidor.  
Om det bara är en enda sida som skall få ett annat sidhuvud, kan du också täcka sidhuvudet med en textram.  
Bakgrunden skall ha pappersfärgen "Vit".  
Information om sidhuvuden och sidfötter i HTML-format  
Några av kommandona för sidhuvuden och sidfötter är också tillgängliga för HTML-dokument.  
Eftersom sådana sidhuvuden och sidfötter inte är gjorda för HTML-definitionen exporteras de som speciella taggar.  
De utvärderas korrekt när en HTML-sida laddas med %PRODUCTNAME.  
Webbläsare visar sidhuvudets eller sidfotens innehåll i form av den text som stod där när HTML-exporten gjordes, medan %PRODUCTNAME fogar in ett fältkommando igen och uppdaterar det vid behov. (Författare och avsändare fogas dock bara in som fältkommando om det är du själv som är författare eller var den som ändrade dokumentet senast.) Sidhuvuden och sidfötter exporteras till HTML-dokument om de aktiverats i läget onlinelayout.  
Definiera olika sidhuvuden  
Ett definierat sidhuvud (och sidfot) gäller för alla sidor som tilldelats sidformatmallen.  
Men ofta kanske du behöver olika sidhuvuden för den första sidan och för jämna och ojämna sidor.  
På de vänstra (jämna) sidorna kan t.ex. namnet på kapitlet stå och på de högra (udda) sidorna namnet på det första underordnade kapitlet.  
Eftersom sidhuvudena är en egenskap från sidformatmallarna måste du definiera olika sidformatmallar och tilldela sidorna dem.  
Det finns redan fördefinierade sidformatmallar för Första sidan, Vänstersida och Högersida, som du kan anpassa efter dina behov.  
Sidformatmallen för vänstersidor kan t.ex. ha olika sidmarginaler för invändig och utvändig marginal, och formatmallen för högersidor har samma marginaler, fast spegelvända.  
Om du inte behöver olika sidhuvuden och sidfötter kan du också välja en spegelvänd sidlayout (i listrutan med samma namn under fliken Sida).  
Bytet mellan jämna och ojämna sidformatmallar och mellan Första sidan och Vänstersida sker automatiskt om du definierar en Nästa formatmall.  
Om du definierar sidformatmallen med nästa formatmall och tilldelar den första sidan den nya sidformatmallen för den första sidan, tilldelar %PRODUCTNAME automatiskt de följande sidorna rätt sidformatmallar.  
Öppna ett nytt tomt textdokument  
Klicka på ikonen Sidformatmallar i Stylist.  
Markera formatmallen Första sidan, som du använder som utgångspunkt för din egen sidformatmall.  
Öppna snabbmenyn och välj Nytt.  
Klicka på fliken Administrera i dialogrutan Sidformatmall.  
Välj "Vänstersida" som Nästa formatmall.  
Välj också "Högersida" som Nästa formatmall för "Vänstersida "och "Vänstersida" som Nästa formatmall för "Högersida ".  
Infoga kapitelinformation i sidhuvud.  
I ett dokuments sidhuvud kan du t.ex. infoga fält som innehåller filnamnet, datum och klockslag och rullande kapitelöverskrifter.  
1.  
Skriv ett längre dokument där du använder styckeformatmallarna "Överskrift 1" för kapitelnamnen.  
2.  
Aktivera sidhuvuden för dokumentet (Infoga - Sidhuvud eller Format - Sida - Sidhuvud).  
3.  
Placera markören i sidhuvudet genom att klicka en gång med musen.  
4.  
Skriv "Kapitel:"  
5.  
Välj Infoga - Fältkommando - Andra.  
6.  
I dialogrutan Fältkommandon klickar du på fliken Dokument och väljer fälttypen Kapitel och formatet Kapitelnamn.  
Om du inte vill citera stycken som är formaterade med Överskrift 1, utan med Överskrift 2, anger du 2 under Nivå.  
7.  
Klicka på Infoga för att infoga kapitelnamnet och stäng dialogrutan.  
Nu visas den önskade kapitelöverskriften automatiskt i sidhuvudet på varje sida i ditt dokument.  
På liknande sätt kan du till exempel infoga sidnummer eller datum.  
Du hittar egna menykommandon till det under Infoga - Fältkommando.  
Där väljer du bland kommandona Datum, Klockslag, Sidnummer, Sidantal, Ämne, Titel och Författare.  
Alla ytterligare fältkommandon väljer du under kommandot Andra.  
Infoga linje under sidhuvud  
Du har dessutom möjlighet att använda ytterligare egenskaper om du öppnar dialogrutan Format - Sida och klickar på fliken Sidhuvud.  
Första gången du definierar ett sidhuvud för dokumentet kan du också göra det under fliken Sidhuvud.  
Markera då rutan Sidhuvud på.  
När du stänger dialogrutan med OK skapas ett sidhuvud som du sedan kan fylla med innehåll i dokumentet.  
Om du klickar på kommandoknappen Fler under fliken Sidhuvud kan du göra fler inställningar av sidhuvudets inramning och bakgrund.  
Du definierar en linje under sidhuvudet genom att klicka på fliken Inramning och där klicka mellan de båda nedre vinkelmarkeringarna i den undre rutan i området Linjeplacering.  
Under den här fliken definierar du även stilen på linjen och avståndet mellan texten i sidhuvudet och linjen.  
Dold text  
Du vill att en viss text bara ska visas och skrivas ut när ett villkor uppfylls.  
Villkoret jämför ett fast värde med innehållet i en variabel eller ett databasfält.  
De möjliga operatorerna finns i listan över operatorer.  
Det finns följande möjligheter:  
Dold text - du väljer kommandot Infoga - Fältkommando - Andra - fliken Funktioner och matar i den dolda texten (t.ex. delar av ett stycke).  
Dolt stycke - du väljer kommandot Infoga - Fältkommando - Andra - fliken Funktioner och matar in det dolda stycket.  
Det går också att dölja ett tomt stycke, t.ex. när ett databasfält inte har något innehåll för den aktuella dataposten.  
Du kan visa dolda stycken på bildskärmen oberoende av villkoret genom att markera kommandot Visa - Dolda stycken.  
Villkorlig text - du väljer kommandot Infoga - Fältkommando - Andra - fliken Funktioner och matar in den villkorliga texten.  
För villkorlig text finns det två textalternativ, det ena alternativet visar och skriver ut texten om villkoret är uppfyllt, och det andra när villkoret inte är uppfyllt.  
Dolt område - du definierar områden via kommandot Infoga - Område.  
Ett område kan innehålla flera stycken.  
Området kan döljas oberoende av ett villkor.  
Så här skriver du text som bara är synlig på bildskärmen och inte skrivs ut  
Du gör så här om du bara vill visa text i ditt dokument på bildskärmen, men inte skriva ut den:  
Rita upp en manuell ram.  
Skriv texten i ramen.  
Välj Format - Ram....  
Du ser dialogrutan Ram.  
Ta bort markeringen framför rutan Skriv ut under fliken Tillägg.  
Ramen visas bara på bildskärmen och skrivs inte ut.  
Infoga - Fältkommando - Andra  
Infoga - Område  
Infoga hyperlänk i textdokument från Navigator  
Infoga hyperlänk med hjälp av Navigator  
Draläget Infoga som hyperlänk måste vara aktiverat.  
På det här sättet kan du också infoga hyperlänkar till objekt i andra öppnade dokument.  
Om du t.ex. vill infoga en hänvisning av typen "se illustration 3" i din text, gör du så här:  
Öppna Navigator  
Klicka på plustecknet bredvid illustrationerna i Navigator  
Välj draläget Infoga som hyperlänk (om det inte redan är markerat)  
Dra posten "Illustration 3" till textdokumentet.  
I textdokumentet infogas namnet på illustrationen som understruken hyperlänk.  
Genom att klicka kan du hoppa direkt till illustrationen.  
Om "Illustration 3", som hyperlänken ska hänvisa till, finns i ett annat textdokument, gör du så här:  
Öppna båda dokumenten  
Öppna Navigator i det textdokument där du vill infoga hyperlänken.  
Välj det andra textdokumentet, som innehåller illustrationen, i kombinationsfältet längst ner i Navigator.  
Välj draläget Infoga som hyperlänk  
Klicka på plustecknet bredvid illustrationerna i Navigator  
Dra posten "Illustration 3" till textdokumentet.  
Importera en punktuppställning från andra ordbehandlingsprogram  
Alla ordbehandlingsprogramm har sina egna sätt att administrera punktuppställningar och numreringar internt.  
Om importfiltret i %PRODUCTNAME inte skulle utvärdera den här informationen korrekt, gör du så här.  
Importera dokumentet från det andra programmet (Arkiv - Öppna - listrutan Filtyp).  
Om punkterna inte importeras korrekt, kan du försöka spara dokumentet i RTF-format i det andra programmet och importera dokumentet igen.  
Markera och kopiera strängen, som nu står i början av varje punktuppställning, till urklippet.  
Det kan t.ex. vara en stjärna * följt av en tabb.  
Öppna dialogrutan Sök och ersätt.  
Klistra in urklippets innehåll i fältet Sök efter.  
Du kan se till att söktexten bara hittas i början av stycken genom att infoga ett ^ framför söktexten och markera rutan Reguljärt uttryck.  
Klicka på Sök alla.  
Nu markeras alla importerade punktuppställningar.  
Stäng inte dialogrutan Sök och ersätt än.  
Klicka på ikonen Punktuppställning på / av på textobjektlisten.  
Nu omvandlas alla importerade punktuppställningar till %PRODUCTNAME -punktuppställningar.  
Klicka på Ersätt alla i dialogrutan Sök och ersätt.  
Eftersom fältet är tomt, raderas alla markerade strängar med t.ex. stjärna * och tabb.  
I dialogrutan Format - Numrering / Punktuppställning kan du definiera typ av punkter för punktuppställningarna.  
Redigera eller radera förteckningspost  
De förteckningsposter som du definierat är markerade med grått i dokumentet för att de skall vara lättare att hitta.  
Markeringarna skrivs inte ut.  
Om du inte heller vill att de ska visas på bildskärmen kan du ta bort dem via Visa - Markeringar.  
Om du vill redigera en post placerar du markören omedelbart framför eller i den aktuella posten.  
Sedan väljer du Redigera - Förteckningspost.  
Du kan ändra texten i textfältet Post.  
Du kan radera den här posten från listan med kommandoknappen Radera.  
Om du ändrar den visade texten i posten kommer den ändrade texten att infogas i den genererade förteckningen.  
På postens ställe i dokumentet visas då bara en smal grå markering.  
Om du vill redigera en sådan post placerar du markören omedelbart bakom markeringen och väljer Redigera - Förteckningspost.  
Med pilknapparna i dialogrutan Redigera förteckningspost växlar du till nästa eller föregående post av samma förteckningstyp.  
Uppdatera, redigera eller radera förteckning  
Placera markören i förteckningen och öppna snabbmenyn.  
På snabbmenyn finns kommandon för att uppdatera, redigera eller radera den aktuella förteckningen.  
Förteckningar är skyddade mot ändringar i förinställningen.  
Du kan bara placera markören i förteckningen om rutan Markör i skyddade områden - Tillåt under Verktyg - Alternativ - Textdokument - Formateringshjälp är markerad.  
Om du vill redigera förteckningen öppnar du snabbmenyn på förteckningen och väljer Redigera förteckning.  
I dialogrutan klickar du på fliken Förteckning och avmarkerar rutan Skyddad mot manuella ändringar.  
Definiera förteckningsposter  
Innan du skapar en förteckning definierar du posterna som ska tas med i förteckningen.  
Det är enklast med poster i en innehållsförteckning: tilldela dina överskrifter styckeformatmallarna "Överskrift 1" till "Överskrift 10 ", beroende på hierarkinivå.  
Innehållsförteckningen kan då skapas automatiskt. (Du kan även lägga till stycken som är formaterade med andra styckeformatmallar i innehållsförteckningen, se.)  
Poster för andra förteckningar definierar du först som poster i dokumentet.  
Markera det eller de ord som skall tas med i förteckningen.  
Du kan hålla ner skifttangenten och markera flera ord om de står efter varandra, eller hålla ner Kommando Ctrl -tangenten när du markerar om orden är utspridda.  
Vid ett enstaka ord räcker det att ställa markören i ordet.  
Ta med de markerade orden i en förteckning med Infoga - Förteckningar - Post.  
I fältet Post anger du det som ska stå i förteckningen.  
Du kan t.ex. skriva "Lexikon, definiera" medan det bara står "Lexikon "i texten.  
Du definierar alla likadana ord i en text som poster om du markerar rutan Använd på alla liknande texter i dialogrutan Infoga - Förteckningar - Post.  
Om du vill ta med orden i en egen förteckning klickar du på ikonen Ny användardefinierad förteckning i dialogrutan Infoga förteckningspost.  
Du ser en dialogruta där du kan ange förteckningens namn.  
Det här namnet blir senare förteckningens rubrik.  
Du kan ändra rubriken för en förteckning utan att innehållet i förteckningen påverkas.  
Redigera förteckningsformat  
I dialogrutan Infoga förteckning kan du även redigera förteckningens format under fliken Poster.  
Här kan du bl.a. ändra hur poster, tabbar och sidnummer är placerade.  
Under fliken Mallar kan du tilldela andra styckeformatmallar.  
Det finns mer information i %PRODUCTNAME -hjälpen.  
Du kan automatiskt tilldela posterna i innehållsförteckningen hyperlänkar.  
Placera sedan markören efter <E> och klicka en gång till på Hyperlänk.  
I dokumentets innehållsförteckning kan du sedan klicka på en hyperlänk för att komma direkt till den första sökträffen.  
För att den här funktionen skall fungera måste innehållsförteckningen vara skapad av överskrifter.  
Skapa sakregister  
Placera markören på stället i texten där sakregistret ska skapas.  
Välj Infoga - Förteckningar - Förteckningar.  
Dialogrutan Infoga förteckning visas.  
Klicka på fliken Förteckning och välj typen "Sakregister".  
Klicka på OK om du vill generera sakregistret med standardinställningarna.  
Du kan t.ex. välja om de bokstäver under vilka poster står skall framhävas som mellanrubriker ("Alfabetiskt skiljetecken "under fliken Poster), eller om det skall göras skillnad mellan stora och små bokstäver och mycket annat.  
Om du vill ändra formateringen av de enskilda raderna i förteckningen är det bäst om du redigerar styckeformatmallarna i Stylist.  
Alla direkta formateringar skrivs över vid nästa uppdatering.  
Använda konkordansfil  
Om du vill kan du lägga till uppslagsord från en konkordansfil.  
I en konkordansfil är ett antal uppslagsord förtecknade och det finns uppgifter om hur de här uppslagsorden ska visas i sakregistret.  
Välj Infoga - Förteckningar - Förteckningar.  
Under fliken Förteckning väljer du typen Sakregister.  
Markera rutan Konkordansfil.  
Genom att klicka på kommandoknappen Fil kan du nu välja om du vill öppna en konkordansfil, skapa en ny eller redigera en konkordansfil.  
Det finns mer information om konkordansfilens struktur i %PRODUCTNAME -hjälpen.  
Skapa litteraturförteckning  
En litteraturförteckningspost kan t.ex. se ut så här i text: "Smith [Smith 1995] har också studerat denna fråga ingående".  
Läsaren vet då att han kan hitta närmare uppgifter (författarens fullständiga namn, boktitel, förlag o.s.v.) i litteraturförteckningen under stickordet [Smith 1995].  
Under fliken Poster i dialogrutan Infoga förteckning (typ "Litteraturförteckning") kan du själv välja vilka uppgifter som ska stå i litteraturförteckningen.  
Du behöver andra uppgifter i t.ex. poster för tidskriftsartiklar än i poster för böcker.  
Därför är litteraturdatabasen indelad i olika typer av litteraturkällor.  
När du vill redigera litteraturdatabasen väljer du Verktyg - Litteraturdatabas.  
Du kan också skapa en datapost i dialogrutan Infoga post i litteraturförteckning (med kommandoknappen Ny).  
De sparas dessutom bara om du verkligen infogar den nya posten.  
Du skapar litteraturförteckningsposterna i texten genom att placera markören där posten ska stå och sedan välja Infoga - Förteckningar - Litteraturförteckningspost.  
Följande dialogruta visas:  
Bestäm först om du vill välja posten från dataposterna i litteraturdatabasen eller från posterna som finns i det aktuella dokumentet (och som kan skilja sig från likalydande poster i litteraturdatabasen).  
En post i dokumentinnehållet kan vara likadan som en post i litteraturdatabasen.  
Posten i dokumentet har högre prioritet.  
Om den önskade posten redan finns som datapost väljer du den i listrutan Kort beteckning och klickar på Infoga.  
Om den önskade posten inte finns än skapar du en ny post.  
Om du använder kommandoknappen Ny kan du definiera en ny datapost, som bara är känd i det aktuella dokumentet.  
Om dataposten ska finnas med i din litteraturdatabas, väljer du Verktyg - Litteraturdatabas, anger den nya dataposten där och infogar sedan litteraturförteckningsposten i dokumentet.  
Förteckning över flera dokument  
Om du vill skapa en förteckning över flera dokument, finns det flera möjligheter:  
Du kan skapa en förteckning i varje enskilt dokument och kopiera förteckningarna till ett dokument och redigera dem.  
Ett ännu bättre sätt är att markera varje enskild förteckning som område (Infoga - Område) och infoga dessa områden som länk i ett gemensamt förteckningsdokument.  
Om du arbetar med ett samlingsdokument kan du skapa gemensamma förteckningar över samtliga deldokument.  
Skapa innehållsförteckning  
Placera markören där innehållsförteckningen ska skapas.  
Välj Infoga - Förteckningar - Förteckningar.  
Dialogrutan Infoga förteckning visas.  
Under fliken Förteckning väljer du typen "Innehållsförteckning" (första gången dialogrutan öppnas är fliken och typen redan förvald).  
Klicka på OK när du vill generera innehållsförteckningen av överskrifterna och de förteckningsmarkeringar som du har definierat.  
Om du vill ta med fler stycken med andra styckeformatmallar i innehållsförteckningen kan du markera fältet Ytterligare mallar och klicka på ikonen efter fältet.  
Då öppnas en dialogruta där du kan definiera för varje styckeformatmall i dokumentet om den ska visas i innehållsförteckningen och på vilken nivå.  
Om du ändrar överskrifterna senare, ändrar deras ordningsföljd eller fogar in nya kapitel måste du uppdatera innehållsförteckningen.  
Placera textmarkören i innehållsförteckningen.  
Öppna snabbmenyn och välj Uppdatera förteckning.  
Du kan också välja Verktyg - Uppdatera - Alla förteckningar för att uppdatera alla förteckningar samtidigt.  
Skapa användardefinierade förteckningar  
Du kan skapa hur många egna förteckningar som helst.  
I dialogrutan Infoga förteckningspost kan du klicka på ikonen Ny användardefinierad förteckning och sedan ange namnet på den nya förteckningen.  
Sedan lägger du till posterna för den nya förteckningen.  
Slutligen kan du skapa förteckningen i ditt dokument:  
Placera markören på det ställe i texten där den användardefinierade förteckningen ska skapas.  
Välj Infoga - Förteckningar - Förteckningar...  
Dialogrutan Infoga förteckning visas.  
Klicka på fliken Förteckning och välj typen "Användardefinierad".  
Om du har gett den egna förteckningen ett namn väljer du namnet i listrutan Typ.  
Klicka på OK när du vill skapa förteckningen av markeringarna för förteckningen som visas i listrutan Typ.  
Välj sedan någon av de mallar som används i dokumentet, om du vill skapa förteckningen av alla stycken som är formaterade med den här mallen.  
Markera de andra rutorna i området Skapa från om du vill skapa förteckningen av alla objekt av en viss typ.  
Ge förteckningen ett passande namn i fältet Rubrik. (Du kan också ändra namnet direkt i dokumentet men då skrivs det över när förteckningen uppdateras nästa gång.)  
I förteckningen visas objektens namn som du har tilldelat objekten under fliken Tillägg i respektive egenskapsdialog.  
Infoga stycke ovanför tabell i början av sidan  
Har du infogat en tabell i början av ett textdokument eller direkt efter en fast sidbrytning och vill nu infoga text framför den här tabellen?  
Placera markören i den första cellen i tabellen, alldeles i början av det eventuella innehållet i den här cellen.  
Tryck på returtangenten där.  
Tabellen flyttas en rad ner.  
Om du vill radera den här raden framför tabellen sätter du textmarkören i den (tomma) raden och trycker på Delete.  
Infoga ett grafikobjekt per dialogruta  
Placera markören på det ställe i dokumentet där du vill infoga grafikobjektet.  
Välj Infoga - Grafik - Från fil.  
Dialogrutan Infoga grafik öppnas.  
Välj ut ett grafikobjekt och klicka på Öppna.  
I standardinställningen infogas grafikobjektet centrerat ovanför det aktuella stycket.  
Infoga ett diagram från %PRODUCTNAME Calc  
Dra och släppa en kopia av ett diagram  
Öppna %PRODUCTNAME Writer-dokumentet där du vill infoga ett diagram.  
Öppna %PRODUCTNAME Calc-dokumentet som innehåller diagrammet.  
Markera diagrammet genom att klicka på det en gång.  
Diagrammet får åtta handtag.  
Om du dubbelklickar på diagrammet av misstag, sätts det i redigeringsläge vilket du kan se på den gråa kanten.  
Klicka en gång utanför diagrammet för att lämna redigeringsläget.  
Dra diagrammet till %PRODUCTNAME Writer-dokumentet.  
Om %PRODUCTNAME Writer-dokumentet inte är synligt direkt, kan du ordna fönstren först.  
Om ditt operativsystem eller din fönsterhanterare har ett aktivitetsfält, kan du först dra diagrammet till kommandoknappen för %PRODUCTNAME Writer-dokumentet på aktivitetsfältet, fortsätta att hålla ner musknappen och vänta där tills %PRODUCTNAME Writer-fönstret öppnas i förgrunden och sedan dra till dokumentet.  
I %PRODUCTNAME Writer-dokumentet placerar du diagrammet eller ändrar storleken, precis som med andra objekt.  
Om du vill ändra data i diagrammet i efterhand, dubbelklickar du på det och redigerar sedan data och andra egenskaper.  
Diagram med länkade data  
Om diagrammet har infogats enligt metoden som beskrivs ovan uppdateras det inte om data ändras i %PRODUCTNAME Calc-dokumentet.  
Om det är viktigt att diagrammet ständigt uppdateras kan du göra så här:  
Kopiera cellområdet, som du vill skapa diagrammet av, från Calc-dokumentet till urklippet.  
Växla till Writer-dokumentet och klicka länge på ikonen Klistra in på funktionslisten.  
På undermenyn väljer du "DDE-länk".  
Uppgifterna finns nu i en texttabell i Writer-dokumentet och är hela tiden länkade till källdata i Calc-dokumentet via DDE.  
Sätt markören i texttabellen i Writer-dokumentet.  
Klicka på ikonen Infoga diagram på utrullningslisten Infoga objekt på verktygslisten.  
Infoga grafik från %PRODUCTNAME Draw eller Impress  
Om du vill infoga ett grafikobjekt från ett dokument i ett annat dokument, kan du kopiera grafikobjektet genom att använda dra-och-släpp.  
Om du vill publicera ditt dokument bör du följa lagen om upphovsrätt och inhämta tillstånd från författarna till originalsidan för säkerhets skull.  
Öppna dokumentet där du vill infoga grafikobjektet.  
Öppna dokumentet som du vill kopiera grafikobjektet från.  
Håll ner Alternativ Alt -tangenten och klicka på grafikobjektet så att det markeras, men utan att en hyperlänk som eventuellt är kopplad till det aktiveras.  
Håll ner musknappen och vänta ett ögonblick medan grafikobjektet kopieras till urklippet.  
Dra grafikobjektet till det andra dokumentet.  
Om dokumenten inte är synliga bredvid varandra, drar du först muspekaren till måldokumentets kommandoknapp.  
Fortsätt att hålla ner musknappen!  
Dokumentet aktiveras och visas och du kan föra muspekaren till dokumentet.  
Släpp musknappen så snart den gråa textmarkören antyder den plats där du vill infoga grafikobjektet.  
En kopia av grafikobjektet infogas.  
Om grafikobjektet är kopplat till en hyperlänk infogas hyperlänken i stället för grafikobjektet.  
Infoga ett grafikobjekt från Gallery med dra-och-släpp  
Dra ett grafikobjekt från Gallery till ett text-, tabell - eller presentationsdokument, så infogas grafikobjektet där.  
Om du släpper grafikobjektet direkt på ett ritobjekt gäller följande:  
Om du drar utan tilläggstangent (det finns inget tilläggstecken vid muspekaren) överförs bara teckenattributen från Gallery och tilldelas ritobjektet på vilket du släpper musknappen.  
Om du håller ner Ctrl-tangenten när du drar (du ser ett plustecken vid muspekaren) infogas grafikobjektet som objekt.  
Om du håller ner Skift+Ctrl-tangenterna (du ser en länkningspil vid muspekaren) ersätts ritobjektet av grafikobjektet från Gallery, men det ersatta ritobjektets position och storlek bibehålls.  
Infoga ett grafikobjekt med skanner  
Förutsättningen för att du ska kunna skanna i %PRODUCTNAME är att du har installerat en skanner med lämpligt drivrutinsprogram i ditt system.  
I Windows understödjer %PRODUCTNAME TWAIN-standarden.  
I Unix understödjer %PRODUCTNAME SANE-standarden.  
Placera markören på det ställe i dokumentet där du vill infoga grafikobjektet.  
Välj Infoga - Grafik - Skanna.  
På undermenyn finns ett kommando som öppnar en dialogruta där du kan välja skanningskälla.  
Välj kommandot som startar skanningen på undermenyn.  
Skanningsdrivrutinen öppnar sitt fönster där du följer skannertillverkarens anvisningar.  
När skanningen är avslutad har bilden infogats i %PRODUCTNAME -dokumentet.  
Infoga grafik  
Det finns flera olika sätt att infoga ett grafikobjekt i ett textdokument:  
Infoga horisontell linje  
Via menykommandot Infoga - Horisontell linje öppnar du en dialogruta där du kan välja linjer.  
Linjerna är grafikobjekt som är förankrade vid det aktuella stycket och som är centrerade mellan sidmarginalerna.  
Linjerna finns också i ett tema i Gallery.  
Om du vill använda en linje från Internet, lägger du till den till motsvarande tema i Gallery.  
Sedan går det att välja linjen i den här dialogrutan.  
Gallery  
Ändra numrering via tangentbordet  
Om du vill flytta en numrering ett steg längre ner (eller flytta den åt höger) i hierarkin placerar du markören i början av det numrerade stycket och trycker på tabbtangenten.  
Med skifttangent plus tabbtangent flyttas en punktuppställning eller numrering med indrag upp ett steg (åt vänster) igen.  
Om du vill infoga en tabb i början av en numrerad rad, använder du Kommando Ctrl +Tabb.  
Slå ihop två separata numreringar  
Om du vill slå ihop två separata numreringar till en genomgående numrering, markerar du båda numreringarna och klickar sedan två gånger efter varandra på ikonen Numrering på / av på objektlisten.  
Exempel  
Sedan har du omvandlat punkt 3 till ett stycke utan numrering.  
Numreringen ser nu ut så här:  
1.  
Första raden  
2.  
Andra raden  
Tredje raden  
1.  
Fjärde raden  
2.  
Femte raden  
Radera den tredje raden helt och hållet så fortsätter numreringen inte automatiskt från 1. till 4..  
Markera raderna som är numrerade med 1., 2., 1., 2. och klicka sedan två gånger efter varandra på ikonen Numrering på / av på objektlisten.  
Placera markör vid bokmärke  
Om det finns bokmärken i ett textdokument, kan du öppna en snabbmeny med dem genom att hålla ner Ctrl-tangenten och klicka med musen klicka med den högra musknappen i fältet Sida på statuslisten.  
Om du klickar på ett av bokmärkena i snabbmenyn flyttar du textmarkören dit.  
Infoga bokmärke  
Definiera linjeslut  
Rita linjeslutet med hjälpmedlen från utrullningslisten Ritfunktioner och lägg till det i listan med linjeslut.  
Rita ett objekt som passar som linjeslut med hjälp av ritfunktionerna.  
Objektets spets ska peka uppåt.  
Öppna dialogrutan Format - Linje medan objektet fortfarande är markerat.  
Välj fliken Linjeslut.  
Klicka på Lägg till.  
Ge det nya slutet ett nytt namn.  
Linjeslutet sparas automatiskt.  
Rita linje i text  
Linjerna kan ha valfri form, bredd och färg och andra attribut.  
En horisontell linje som är lämplig för webbsidor skapar du genom att tilldela ett tomt stycke det medföljande styckeformatet Horisontell linje.  
Placera markören i det tomma stycket och dubbelklicka sedan på Horisontell linje i Stylist.  
Om du inte hittar den bland styckeformaten i Stylist kan du välja "Alla mallar" i stället för "Automatiskt ".  
En linje direkt ovanför, bredvid eller under ett stycke ritar du med Format - Stycke - Inramning.  
Den här funktionen förklaras utförligt i %PRODUCTNAME -hjälpen.  
Men om du vill definiera attributen och riktningen för en linje själv, så använder du ritobjektet Linje på följande sätt:  
1.  
Öppna utrullningslisten Visa ritfunktioner på verktygslisten och klicka på ikonen Linje.  
Muspekaren blir till ett hårkors med en linje.  
2.  
Klicka på startpunkten för linjen i dokumentet, håll ner musknappen och dra tills du har nått slutpunkten för linjen.  
Om du håller ner skifttangenten samtidigt, kan du bara rita horisontella, vertikala och diagonala linjer.  
3.  
Släpp musknappen när linjen har den riktning och längd som du vill ha.  
Du kan rita fler linjer direkt.  
Avsluta funktionen via Esc-tangenten eller genom att klicka på ikonen Urval på utrullningslisten Visa ritfunktioner.  
4.  
När du har klickat på ikonen Urval kan du hålla ner skifttangenten och markera alla linjer samtidigt för att sedan till exempel tilldela dem en färg, bredd eller andra attribut.  
De kan i stället exporteras som grafik.  
Format - Stycke - Inramning  
Definiera linjestil  
Markera ett ritobjekt som du t.ex. har ritat med hjälp av utrullningslisten Visa ritfunktioner.  
Öppna dialogrutan Format - Linje.  
Klicka på fliken Linjestil.  
Här definierar du en linjestil.  
Som du ser finns det många olika möjligheter att kombinera streck, punkter och avstånd.  
Punkter är alltid lika långa som breda, medan du fritt kan ställa in längden på streck och avstånd.  
Om du markerar rutan Anpassa till linjebredd kan du ställa in längderna i procent av linjebredden.  
Definiera en ny linjestil och klicka på Lägg till.  
Ge den nya stilen ett namn.  
Den nya stilen sparas automatiskt.  
Du kan spara linjestilen i en egen linjestilstabell.  
Om du öppnar dialogrutan Spara som via symbolen Spara linjestiltabell, sparas alla tillgängliga linjestilar som fil med ett namn som du väljer.  
Använd linjestilar  
Markera det objekt som du vill tilldela en ny linjestil.  
Öppna till exempel utrullningslisten Ritfunktioner och rita en linje.  
Linjen är markerad när du har ritat den.  
Nu kan du tilldela linjen attribut på olika sätt.  
I ritobjektlisten hittar du ikoner och listrutor för att välja olika attribut.  
I snabbmenyn och i menyn Format kan du välja kommandot Linje.  
På ritobjektlisten kan du öppna dialogrutan Format - Linje... genom att klicka på ikonen Linje.  
Om du klickar på den får du i en utrullningslist se ett urval av de tillgängliga linjesluten för höger och vänster.  
Klicka på de önskade symbolerna.  
Själva linjestilen väljer du i listrutan Linjestil och bredden med rotationsknapparna för Linjebredd.  
Om det står 0,00 cm här, visas linjen med en bredd på 1 pixel.  
I nästa listruta Linjefärg väljer du färg för linje och linjeslut.  
Om du öppnar dialogrutan Linje kan du göra önskade inställningar under flikarna.  
Du kan också ladda linjestil - och linjesluttabeller med olika stilar och ändar.  
De olika alternativen beskrivs utförligt i %PRODUCTNAME -hjälpen.  
Sätta på och stänga av hyperlänk  
Håll ner Alternativtangenten Alt-tangenten och klicka på hyperlänken.  
På statuslisten för textdokument finns fältet HYP eller SEL.  
Du kan växla mellan HYP och SEL genom att klicka i fältet.  
När HYP visas, utförs en hyperlänk när du klickar på den.  
Om SEL visas, kan du klicka på hyperlänken och redigera den.  
Du trycker in ikonen Utkastläge på / av på utrullningslisten Formulärfunktioner.  
Kopiera formatmallar i dokument  
Du kan ladda formatmallarna från ett annat dokument i det aktuella dokumentet.  
Välj Format - Mallar - Ladda och välj ett dokument.  
Välj om du vill överföra textformatmallar (det är styckeformatmallar och teckenformatmallar), ramformatmallar, sidformatmallar och / eller numreringsformatmallar och om mallarna i det aktuella dokumentet ska skrivas över av de nya mallarna.  
Om du klickar på kommandoknappen Från fil... öppnas en dialogruta där du kan välja mall på samma sätt som under Arkiv - Nytt - Mallar och dokument.  
Skapa standardbrev  
Här följer en snabb och en utförlig beskrivning av hur standardbrev (kopplad utskrift) skapas:  
Snabb beskrivning (för snabbt resultat)  
Registrera en adressdatakälla i %PRODUCTNAME om du inte redan har gjort det.  
Det finns en beskrivning under sökordet Adressbok i %PRODUCTNAME -hjälpen.  
Öppna en av mallarna för standardbrev (kopplad utskrift) med Skift+Ctrl+N.  
Mallen Klassiskt brev i kategorin Affärskorrespondens är lämplig.  
Välj ut eller mata in adresserna som ska användas till standardbrevet.  
Låt %PRODUCTNAME skapa och skriva ut standardbreven med kopplad utskrift.  
Utförlig beskrivning (med bakgrundsinformation)  
Till ett standardbrev behöver du dels mottagarnas adresser, som bör vara i form av en databastabell, dels ett textdokument.  
Det står fältkommandon på de ställen i texten där adressen och tilltalet skall skrivas ut i standardbrevet.  
Fältkommandona refererar till motsvarande databasfält och kan definieras i dialogrutan Fältkommando som du öppnar med Infoga - Fältkommando - Andra....  
Fältkommandon är en typ av platshållare i ditt dokument.  
De kan antingen fyllas med aktuella data första gången fältkommandot infogas eller när dokumentet öppnas eller skrivs ut.  
Du kan även utföra en uppdatering för hand, t.ex. med tangenten F9.  
Fasta och variabla fältkommandon  
Fältkommandon som bara fylls med innehåll en gång, nämligen när fältkommandot infogas i dokumentet, är "fasta" fält.  
Du använder t.ex. ett fast datum om du skriver en faktura som baserar på en fakturamall.  
I samma ögonblick som du skapar fakturadokumentet, infogas det aktuella datumet där fältkommandot är placerat och ändras sedan inte mer, eftersom fakturadatumet redan är definierat.  
Ett variabelt datum uppdateras däremot varje gång dokumentet öppnas och skrivs ut.  
Om du uppdaterar fältkommandon för hand, t.ex. med funktionstangenten F9, ställs ett datum in som infogades som fältkommando "variabelt datum" för den aktuella dagen.  
Om du t.ex. vill infoga ett datum som fältkommando i ditt standardbrev, måste du bestämma om det skall infogas som fast eller variabelt fältkommando:  
Välj det fasta datumet om det inte skall ändras igen, alltså om du hade kunnat skriva datumet som klartext (utan fältkommando).  
Vad är fördelen med fältkommandon?  
Du kan spara standardbrevet som dokumentmall senare och om du definierar ett nytt standardbrev som baserar på den här dokumentmallen vid en ännu senare tidpunkt, har du redan automatiskt aktuellt dagsdatum i det nya standardbrevet.  
Om du väljer det variabla datumet som fältkommando, sätts aktuellt datum in varje gång dokumentet öppnas och skrivs ut.  
Förutom datum finns det ett stort antal andra fältkommandon som du kan ha mycket användning för i standardbrev.  
De viktigaste fältkommandona är naturligtvis de som definierar var i brevet vilka delar av mottagaradressen skall infogas.  
De här fältkommandona skapar en direkt förbindelse till databastabellen som innehåller dina mottagaradresser.  
För varje önskat datafält (t.ex. LASTNAME, ADDRESS, CITY) infogas ett eget fältkommando i standardbrevdokumentet.  
När dokumentet skrivs ut sätter %PRODUCTNAME Writer in de önskade datafälten i fältkommandona för varje datapost.  
Om du vill skapa ett helt nytt dokument som innehåller fältkommandona för standardbrev, kan du göra det med dra-och-släpp:  
Öppna textdokumentet och visa den önskade databastabellen med F4.  
Nu kan du peka med musen på ett kolumnhuvud och dra det med nertryckt musknapp till dokumentet.  
Fältkommandot som används till att infoga det här fältet från databastabellen placeras ut automatiskt.  
Välj Arkiv - Nytt - Mallar och dokument och öppna ett dokument som baserar på dokumentmallen Klassiskt brev i kategorin Affärskorrespondens.  
Ett standardbrev som baserar på dokumentmallen "Klassiskt brev" visas.  
Det innehåller redan flera fältkommandon för adress, datum, avsändare och så vidare.  
Dialogrutan Användning av den här mallen visas automatiskt.  
Välj alternativet Flera mottagare (adressdatabas).  
Eftersom adressdatabasen redan är länkad till dokumentmallen "Klassiskt brev", har adresstabellen öppnats automatiskt i datakällvyn.  
Om det inte skulle vara så, kan du öppna datakällan till det aktuella dokumentet genom att trycka på F4.  
Markera dataposterna för vilka du vill skriva ut standardbrev i området med radhuvuden.  
Du kan använda tangenterna Skift och / eller Kommando Ctrl när du klickar, precis som när du markerar i andra listor.  
Om du vill skriva ut standardbrev för alla dataposter i tabellen, klickar du bara på det lilla fältet utan text ovanför radhuvudena.  
Klicka nu på ikonen Kopplad utskrift på databaslisten uppe i datakällvyn.  
Du ser dialogrutan Kopplad utskrift där du väljer vad du vill skicka till skrivaren eller som e-brev.  
Här kan du välja igen om du vill skriva ut de markerade dataposterna, alla dataposter eller ett visst område.  
Om du vill skriva ut ett visst område, t.ex. dataposterna nummer 1 till 5, bör du se till att numren motsvarar ordningsföljden som visas i datakällvyn.  
Vid behov kan du sortera eller filtrera dataposterna i datakällvyn genom att klicka på ikonerna på databaslisten.  
Placera markören i ett datafält som du vill använda till sortering.  
För att till exempel sortera alla dataposter efter postnummer, placerar du markören i en valfri datapost i datafältet POSTALCODE och sedan klickar du på ikonen Sortera stigande.  
Nu är standardbrevet färdigt.  
Avancerade standardbrevfunktioner  
Undvika tomma stycken  
Om du har valt COMPANY som fält för kopplad utskrift i ditt mottagarfält, kan det hända att raden är tom vid utskrift.  
Det sker om databasfältet COMPANY är tomt i databasen.  
Men det går att undvika de här tomma styckena.  
Placera markören framför fältet för kopplad utskrift, COMPANY, i ditt textdokument.  
Öppna dialogrutan Fältkommandon.  
Klicka på fliken Funktioner och välj fälttypen Dolt stycke.  
För nu in följande text i fältet Villkor (utan citationstecken)  
not( COMPANY)  
Om databasfältet COMPANY nu är tomt, skrivs inte raden COMPANY ut, och de resterande fälten flyttas en rad uppåt.  
Arkiv - Kopplad utskrift  
Anvisningar för %PRODUCTNAME Writer  
Mata in och formatera texter  
Mata in och formatera texter automatiskt  
Använda formatmallar, numrera sidor, fältkommandon  
Redigera tabeller i texter  
Bilder, teckningar, clip art, FontWork  
Innehållsförteckning, sakregister  
Överskrifter, numreringar  
Sidhuvuden, sidfötter, fotnoter  
Redigera andra objekt i texter  
Rättstavning, ordlistor, avstavning  
Standardbrev (kopplad utskrift), etiketter och visitkort  
Arbeta med dokument  
Övrigt  
Navigator för textdokument  
Hur kan man visa en översikt där man kan se de olika objekten (t.ex. grafiker eller tabeller) i textdokument?  
Med hjälp av Navigator (F5) kan du få fram en översikt över texten.  
I dokumentet kan du enkelt navigera mellan de olika objekten (stycken, grafiker, tabeller osv.) genom att dubbelklicka på respektive post i Navigator.  
Navigator  
Stänga av taligenkänning i tabell  
Om du matar in ett tal i en texttabell, kan %PRODUCTNAME Writer omvandla talet till ett datum automatiskt.  
Datumformatet, som är definierat i operativsystemet, bestämmer vilket tecken som leder till en automatisk ersättning och hur den formateras.  
I USA används snedstreck som datumavgränsare.  
Om du matar in talet 2 / 28 i ett %PRODUCTNAME Writer i ett amerikanskt operativsystem, omvandlas det här talet automatiskt till datumet 2 / 28 / 01 (år 2001).  
I Tyskland används punkt som datumavgränsare.  
Om du matar in talet 28.2 i %PRODUCTNAME Writer i ett tyskt operativsystem, omvandlas det här talet automatiskt till datumet 28.02.01 (år 2001).  
Du kan sätta på och stänga av ersättningen på följande sätt:  
Placera markören i en texttabell.  
Klicka på kommandot Taligenkänning.  
Om det finns en bock framför kommandot är taligenkänningen och därmed den automatiska ersättningen aktiverad.  
Alternativt kan du göra så här:  
Välj kommandot Verktyg - Alternativ.  
Klicka på Textdokument - Tabell.  
Markera fälten Taligenkänning och Talformatsigenkänning så aktiveras den automatiska ersättningen.  
Verktyg - Alternativ - Textdokument - Tabell  
Numrera rader  
Du bestämmer egenskaperna för radnumreringen under Verktyg - Radnumrering.  
Med radnumreringen kan du förse raderna i ett dokument med nummer.  
Du kan definiera för hela dokumentet om tomma rader och om rader i textramar ska räknas.  
Du kan bestämma med vilka intervall en numrering ska göras och infoga avgränsare för identifiering av ett visst radnummer mellan de här intervallerna.  
Radnumreringarna visas på bildskärmen och skrivs ut.  
Du kan göra fler inställningar för radnumrering i stycket (Format - Stycke - Numrering) eller i styckeformatmallen.  
Den här möjligheten garanterar ytterligare flexibilitet, eftersom du kan utesluta ett stycke från radnumreringen eller börja om numreringen vid ett stycke med ett valfritt startvärde.  
Radnumrering för alla stycken  
Välj Verktyg - Radnumrering.  
Markera rutan Numrering på.  
Nu numreras alla stycken i dokumentet.  
Radnumrering bara för några stycken  
Aktivera radnumreringen för alla stycken, som beskrivet ovan.  
Öppna Stylist och klicka en gång på styckeformatmallen Standard.  
Öppna snabbmenyn genom att klicka med högra musknappen och välj Ändra.  
Dialogrutan Styckeformatmall: Standard  
Klicka på fliken Numrering.  
Ta bort markeringen framför Räkna med raderna i det här stycket.  
Eftersom alla styckeformatmallar bygger på Standard numreras inget stycke nu (om inte en underordnad styckeformatmall har ändrats).  
Markera alla stycken som ska numreras i dokumentet.  
Välj Format - Stycke - Numrering, markera rutan Räkna med raderna i det här stycket och klicka på OK.  
Verktyg - Radnumrering  
Avbryta och fortsätta numrering  
I en rad automatiskt numrerade stycken ska ett stycke inte ha något nummer, som i följande exempel:  
1. första stycket.  
2. andra stycket.  
Ett stycke utan nummer.  
3. stycke nummer tre.  
Du kan välja bland följande metoder:  
Radera automatisk numrering  
Markera styckena 1 till 4 och klicka på ikonen Numrering på / av.  
Placera markören framför det första tecknet i det tredje stycket.  
Radera ett tecken åt vänster med backstegstangenten.  
Stycket är fortfarande indraget men har inte kvar sitt nummer.  
Det fjärde stycket blir nummer 3.  
Den här metoden leder till att utseendet inte ändras när dokumentet sparas i HTML-format.  
Formatering av stycket  
Markera styckena 1 till 4 och klicka på ikonen Numrering på / av.  
Placera markören i det tredje stycket.  
Klicka på ikonen Numrering på / av igen.  
Det tredje stycket har inte kvar sitt nummer och är inte indraget.  
I HTML-format uppstår två oberoende numrerade listor p.g.a. avbrottet.  
Fortsätta numrering med nytt startvärde  
Numrera styckena 1 till 2 med ikonen Numrering på / av.  
Placera markören i det fjärde stycket.  
Välj Format - Numrering / Punktuppställning och klicka på fliken Alternativ.  
Välj posten "1, 2, 3..." i kombinationsfältet Numrering.  
Välj startvärdet i rotationsfältet Börja med - i det här exemplet är det 3.  
Klicka på OK.  
Definiera nummersekvenser  
Om du vill numrera flera element som hör ihop i ett textdokument, till exempel alla kommentarer, alla varningsmeddelanden, alla citat o.s.v., kan du definiera en egen nummersekvens för varje grupp.  
Exempel  
Skriv texten "Citat nummer" framför det första citatet.  
Välj Infoga - Fältkommando - Andra....  
Välj fälttypen "Nummersekvens" under fliken Variabler.  
Skriv det nya namnet "Citat" under Namn.  
Klicka på Infoga och stäng dialogrutan.  
Nu har du definierat en ny nummersekvens, "Citat", med vilken du kan räkna alla citat automatiskt.  
I fältet Värde kan du definiera ett nytt startvärde för hela nummersekvensen.  
Det kan t.ex. vara praktiskt om det rör sig om ett dokument i en serie av sammanhörande dokument.  
Dina nummersekvenser och bildtexter kan även börja om för varje kapitel.  
I dialogrutorna Infoga bildtext och Fältkommando hittar du en urvalslista där du kan välja på vilken kapitelnivå numreringen ska börja om.  
Infoga och radera sidbrytning  
Infoga sidbrytning  
Placera markören på det ställe där den nya sidan ska börja.  
Tryck på Ctrl+Retur.  
En fast sidbrytning infogas och markören står i början av den nya sidan.  
Radera sidbrytning  
Placera markören framför det första tecknet i det första stycket som kommer efter den fasta sidbrytningen.  
Tryck på Delete.  
Den fasta sidbrytningen raderas.  
Radera sidbrytning framför en texttabell  
Placera markören i tabellen och öppna snabbmenyn.  
Välj kommandot Tabell.  
Dialogrutan Tabellformat öppnas.  
Klicka på fliken Textflöde.  
Dialogrutan Infoga brytning  
Sidformatmall och sidnummer  
Du vill först ha en titelsida utan sidnummer i ett textdokument, sedan flera sidor till innehållsförteckningen med små bokstäver som sidnummer (hur lång innehållsförteckningen kommer att bli vet du inte än) och först sedan kommer sidan 1 med siffror som numrering.  
Arbeta med olika sidformatmallar.  
Olika sidformatmallar är motsvarigheten i %PRODUCTNAME Writer till "avsnittsbrytningar" i andra textprogram.  
Det är bäst att placera sidnumren i sidfötter eller sidhuvuden, inte i den löpande texten, så att sidnumrens position inte ändras när text infogas och raderas.  
Gör på följande sätt:  
Skapa nya sidformatmallar  
Tilldela sidorna sidformatmallar  
Redigera sidformatmallar  
Formatera sidnumren i styckeformatmallen för sidfoten om du vill.  
Skapa sidformatmallar  
1.  
Ladda dokumentet som du vill ange eller ändra sidnummer för.  
Du kan också börja med ett helt nytt textdokument, men då bör du först fylla några sidor med text och göra några sidbrytningar, så att du kan tillämpa arbetssättet som beskrivs här.  
2.  
Öppna Stylist.  
3.  
Välj vyn sidformatmallar i Stylist.  
4.  
Öppna snabbmenyn till en av sidformatmallarna och välj Nytt...  
Du ser dialogrutan Sidformatmall med fliken Administrera.  
Markören står i textfältet Namn och du kan ange namnet på den första nya sidformatmallen direkt.  
5.  
Ange Titelsida och tryck på returtangenten.  
Egenskaperna för de nya sidformatmallarna ändrar du senare.  
6.  
I Stylist väljer du nu Nytt... igen via snabbmenyn och definierar en sidformatmall med namnet Innehållsförteckning.  
7.  
Upprepa samma procedur en tredje gång för den nya sidformatmallen Huvudtext.  
De här namnen är naturligtvis bara exempel - du kan använda vilka namn du vill.  
Nu har du skapat tre nya mallar.  
Tilldela sidformatmall  
1.  
Dubbelklicka på Titelsida i Stylist.  
Därmed har du tilldelat den första sidan den här sidformatmallen.  
Som en bekräftelse på detta ser du namnet Titelsida i fältet Sidformatmall nere i statuslisten.  
Du kan också tilldela sidformatmallar som redan finns via snabbmenyn till fältet Sidformatmall i statuslisten och öppna dem för redigering genom att dubbelklicka med musen.  
När du bläddrar vidare i dokumentet kommer du eventuellt att märka att sidformatmallen Titelsida nu gäller för alla sidor i dokumentet.  
Om t.ex. alla sidor hade sidformatmallen Standard innan, har alla sidor nu den nya mallen efter tilldelningen av en ny sidformatmall.  
Sidformatmallar gäller alltid för alla intilliggande föregående och följande sidor i båda riktningar, tills du gör en sidbrytning med byte av sidformatmall i ditt dokument.  
Om du för in en Nästa formatmall till en sidformatmall under fliken Administrera, bestämmer du att nästa formatmall gäller som sidformatmall efter en sidbrytning (oberoende av om du gör den manuellt eller om den görs automatiskt).  
Du kan alltså välja Innehållsförteckning som nästa formatmall till sidformatmallen Titelsida i exemplet som beskrivs här.  
Då får nästa sida efter titelsidan i varje fall sidformatmallen Innehållsförteckning.  
I det här fallet behöver du inte göra detta via dialogrutan Manuell brytning som beskrivs nedan.  
Men du bör bara välja Innehållsförteckning som nästa formatmall till sidformatmallen Innehållsförteckning, eftersom du inte kan veta i förväg hur många sidor innehållsförteckningen kommer att ha.  
2.  
Placera nu markören i början av sidan där innehållsförteckningen ska börja.  
Här ska du ange en manuell brytning med byte av sidformatmall.  
3.  
Välj Infoga - Manuell brytning.  
Dialogrutan Infoga brytning öppnas.  
4.  
Välj alternativet Sidbrytning som Typ.  
I listrutan väljer du sidformatmallen Innehållsförteckning som skall gälla från och med här.  
Klicka på OK.  
5.  
Placera markören i början av den första raden i huvudtexten.  
6.  
Välj också här Infoga - Manuell brytning....  
Dialogrutan Infoga brytning öppnas.  
7.  
Välj alternativet Sidbrytning som Typ.  
I kombinationsfältet väljer du sidformatmallen Huvudtext som skall gälla från och med här.  
Markera Ändra sidnummer och välj det nya sidnumret 1.  
Klicka på OK.  
Om du vill att sidhuvudena eller sidfötterna ska ha olika innehåll på vänster - och högersidor, räcker det att avmarkera Samma innehåll till höger / vänster.  
Under Format - Sida - Sida kan du välja sidlayouten "Spegelvänt".  
Då kan du bl.a. definiera en inre och yttre marginal för texten.  
Ofta har höger - och vänstersidorna i huvudtexten olika sidformatmallar så att t.ex. vänstersidorna har ett sidhuvud men inte högersidorna.  
Du kan använda dem i stället för Huvudtext.  
Den första sidan i din huvudtext är sida 1 och innehåller formatmallen Högersida.  
Tilldela sedan sidformatmallen Vänstersida som nästa formatmall till Högersida och tvärtom.  
Högersida där du väljer Ändra....  
Under fliken Administrera väljer du nästa formatmall.  
Redigera sidformatmall  
Så här gör du:  
I Stylist väljer du posten Huvudtext, öppnar snabbmenyn och väljer Ändra...  
Dialogrutan Sidformatmall: Huvudtext  
Klicka på fliken Sidfot.  
Klicka på OK.  
Nu ser du en tom sidfot på sidan i ditt dokument.  
Du kan placera markören där genom att klicka med musen.  
När markören står i sidfoten, väljer du Infoga - Fältkommando - Sidnummer.  
Du ser sidnumren som visas i grått på bildskärmen eftersom det är ett fältkommando.  
Om du vill att texten "Sida" skall stå framför sidnumret, placerar du markören framför fältkommandot och matar in texten.  
Klicka på ikonen Centrerat på objektlisten för att centrera det aktuella stycket.  
Sidbrytning som styckeformat  
Att texten automatiskt ska börja med det nya sidnumret 1 har automatiskt förts in som direkt styckeformatering i huvudtextens första stycke.  
Det gäller även om det ännu inte står någon text på den nya sidan efter den manuella brytningen.  
För att kontrollera detta kan du öppna snabbmenyn till det första stycket efter den manuella brytningen och välja Stycke (inte Redigera styckeformatmall eftersom det rör sig om ett direkt formateringsattribut till exakt det här ena stycket).  
Du anger den här egenskapen under Format - Stycke under fliken Textflöde.  
Ändra format på sidnummer  
Även formatet på sidnummer kan du bestämma direkt eller indirekt (som egenskap för sidformatmall) precis som andra textattribut.  
Den direkta formateringen bör du bara använda i undantagsfall.  
Du redigerar ett fältkommando direkt vid den direkta formateringen:  
1.  
Dubbelklicka på fältkommandot med sidnumret.  
Du ser dialogrutan Redigera fältkommando: Dokument  
2.  
Välj formateringen för fältkommandot.  
Klicka på OK.  
Men normalt definierar du formateringen av sidnumren som egenskap till en sidformatmall:  
Öppna snabbmenyn på sidan och välj kommandot Sida.  
Du ser då t.ex. dialogrutan Sidformatmall: Standard  
I stället för "Standard" står namnet på den aktuella sidformatmallen i dialogrutans rubrikrad.  
Klicka på fliken Sida.  
I kombinationsfältet Numrering definierar du hur numreringen skall se ut på alla sidor med den här formatmallen.  
Stäng sedan dialogrutan med OK.  
Nu väljer du formatet Som sidformatmall för fältkommandot som visar sidnumret (se föregående beskrivning av den direkta formateringen).  
Om du vill ändra fler av sidfotens egenskaper, t.ex. teckensnittet, bör du redigera styckeformatmallen Sidfot så att ändringen gäller för alla sidfötter:  
Placera markören i sidfoten.  
Öppna snabbmenyn och välj Redigera styckeformatmall.  
Om du vill öka sidfotens avstånd till texten så är det ett formatattribut i sidformatmallen.  
Ändra sidformatmallen i Stylist via sidformatmallens snabbmeny där du väljer Ändra...  
I dialogrutan Sidformatmall kan du ställa in sidfotens avstånd och höjd.  
Använd inte korrigeringsvärdet som finns under fliken Dokument i dialogrutan "Fältkommandon" som du öppnar via Infoga - Fältkommando - Andra för att ändra sidnumret på en sida.  
Det här värdet är bara till för att t.ex. visa numret på följande sida i slutet av en sida, alltså bara för korrigering av visningen och inte för ändring av själva sidnumret.  
Sidnumret som du har bestämt på en sida (till skillnad från automatiskt satta sidnummer) är en egenskap för den aktuella sidan.  
Egenskapen definieras som direkt formatering vid första stycket på den här sidan.  
Textflöde  
Skapa sidformat liggande  
Öppna Stylist, t.ex. med F11.  
Byt till visningen av Sidformatmallar genom att klicka på ikonen med samma namn.  
Den aktuella sidformatmallen är markerad.  
Klicka på ikonen Ny formatmall från markering.  
Dialogrutan Skapa formatmall visas.  
Ge mallen ett namn.  
Välj t.ex. namnet Liggande och klicka på OK.  
Klicka en gång på den nya mallen Liggande i Stylist.  
Öppna sedan snabbmenyn och välj kommandot Ändra.  
Dialogrutan Sidformatmall: Liggande  
Klicka på fliken Sida, välj alternativet Liggande i området Pappersformat och klicka på OK.  
Nu har du en ny sidformatmall med liggande format som du kan använda på markerade sidor.  
Byta sidformaten stående / liggande  
Du har t.ex. ett 10 sidor långt dokument i stående format, med sidformatet Standard.  
På sidan 5 behöver du liggande format för att få bättre plats med en tabell.  
Skapa en sidformatmall i liggande format.  
Ge den t.ex. namnet Liggande.  
Placera markören direkt framför texten som ska skrivas ut i liggande format.  
Välj kommandot Infoga - Manuell brytning.  
Dialogrutan Infoga brytning.  
Välj alternativet Sidbrytning.  
I kombinationsfältet väljer du sidformatmallen Liggande.  
Klicka på OK.  
Nu har sidorna 1 till 4 standardformat och 5 till slutet av dokumentet liggande format.  
Du placerar alltså markören i slutet av sidan 5 och matar där in en manuell brytning:  
I slutet av sidan med liggande format väljer du kommandot Infoga - Manuell brytning.  
Välj alternativet Sidbrytning.  
I kombinationsfältet väljer du sidformatmallen Standard.  
Klicka på OK.  
I förhandsvisningen kan du kontrollera resultatet: meny Arkiv - Förhandsgranskning / sidutskrift.  
Snabb formatering med intilliggande styckeformat  
Om du har två stycken som kommer efter varandra med olika styckeformat och vill formatera båda samtidigt så går det snabbast om du gör så här:  
Radera styckeslutstecknet mellan de båda styckena.  
Tryck på returtangenten.  
Båda styckena har nu samma format med samma formatmall.  
Om du går till slutet av det första stycket för att radera och trycker på Delete-tangenten där, dras det andra stycket ihop med det första stycket ("Radera åt höger").  
Det andra stycket övertar det första styckets format när du skapar två stycken igen genom att trycka på returtangenten.  
Om du går till början av det andra stycket för att radera och trycker på backstegstangenten (ovanför returtangenten), fixeras det andra stycket ("Radera till vänster"), och när du har tryckt på returtangenten har du två stycken med formatet från det andra stycket.  
Välja pappersmagasin  
Så här kan du välja olika pappersmagasin för dina brev.  
Den första sidan skrivs t.ex. ut med papper från standard-pappersmagasinet där ditt företags brevpapper med fÃ¶retagsbrevhuvud ligger.  
Följande sida skall skrivas ut med papper från pappersmagasin 2 där blankt papper ligger.  
Du tilldelar den första sidan en sidformatmall (i Stylist) och definierar en nästa formatmall till den (under fliken Administrera).  
I egenskaperna för den mallen, under registerflik Sida, har du angivit att papperet skall hämtas från fack 2.  
Om din text blir längre än en sida, använder %PRODUCTNAME automatiskt sidformatmallen som är definierad som nästa formatmall för de följande sidorna.  
Vid utskrift hämtas papperet automatiskt från korrekt pappersmagasin.  
Skriva ut HTML-dokument utan sidhuvud  
Så kan du skriva ut ett HTML-dokument utan sidhuvud / sidfot.  
En dokumentmall används för formatering av HTML-sidor.  
Om du inte vill att sidhuvuden och sidfötter ska skrivas ut när du skriver ut HTML-sidor, måste du ändra den aktuella formatmallen.  
Den heter Standardmall för HTML-filer (html.stw).  
Skapa en säkerhetskopia av filen.  
Öppna dokumentmallen genom att välja filtypen "%PRODUCTNAME %PRODUCTVERSION textdokument" i dialogrutan Öppna.  
Ta bort markeringen i rutan Sidhuvud på.  
%PRODUCTNAME varnar dig nu eftersom du är på väg att kasta bort innehållet i sidhuvudet.  
Bekräfta meddelandet.  
Avslutningsvis klickar du på OK för att stänga sidformat-dialogen.  
Du får då frågan om du vill spara ändringarna.  
När du har gjort detta innehåller HTML-sidor som skrivs ut inga sidhuvuden eller sidfötter längre.  
Förhandsvisning av utskrift  
Innan du skriver ut ett textdokument kan du titta på en förhandsvisning av utskriften så att du t.ex. kan anpassa marginalbredd eller optimera sidbrytningar.  
1.  
Växla till dokumentet som du vill förhandsgranska.  
2.  
Välj Arkiv - Förhandsgranskning / sidutskrift.  
3.  
Anpassa skalan för vyn med hjälp av ikonerna på objektlisten.  
4.  
Bläddra i dokumentet med hjälp av piltangenterna eller ikonerna på objektlisten och kontrollera utskriften.  
Arkiv - Förhandsgranskning / sidutskrift.  
Skriva ut dokument i förminskat format  
Om du vill skriva ut ett textdokument i förminskat format för att spara papper väljer du Arkiv - Förhandsgranskning / sidutskrift.  
Där kan du ställa in om du vill ha två, fyra eller ett valfritt antal dokumentsidor per utskrivet papper bredvid och över varandra.  
Så här skriver du ut två sidor bredvid varandra på ett papper  
1.  
Välj Arkiv - Förhandsgranskning / sidutskrift.  
2.  
I förhandsgranskningen visas två sidor bredvid varandra.  
Om fler eller färre sidor visas klickar du på ikonen Förhandsgranskning: två sidor på objektlisten.  
3.  
Klicka på ikonen Skriv ut förhandsgranskning.  
Bekräfta utskriftsdialogrutan med OK.  
4.  
Om du klickar på ikonen Utskriftsalternativ förhandsgranskning öppnas en dialogruta där du kan göra inställningar för förminskad utskrift.  
Arkiv - Förhandsgranskning / sidutskrift  
Sätta referenser  
Med hjälp av referenser kan du - i motsats till hyperlänkar - bara hänvisa inom samma dokument, inte till andra dokument.  
Referenser anges som fältkommandon.  
Först måste du sätta referensen, d.v.s. definiera målet för en korshänvisning.  
Du kan också sätta korshänvisningar till bildtexter för grafik och tabeller.  
En beskrivning av arbetsstegen följer längre ned.  
Placera markören på det ställe som du vill hänvisa till.  
Markera där ett ord som mål för referensen.  
Det gör det lättare att senare hitta målet för hoppet i dokumentet igen.  
Välj kommandot Infoga - Korshänvisning.  
Välj fälttypen "Sätt referens" och skriv ett entydigt namn för referensen i fältet Namn.  
Klicka på Infoga.  
Nu går du till det ställe där du vill att korshänvisningen ska sättas in.  
Därefter infogar du fältkommandot.  
Välj Infoga - Korshänvisning.  
Välj den här gången fälttypen "Infoga referens".  
I listrutan Urval ser du alla definierade referenser i dokumentet med sina namn.  
Välj önskad referens och ett format och klicka på Infoga.  
Om du vill sätta en referens till ett grafikobjekt eller tabell i det aktuella dokumentet, måste du först infoga en bildtext för grafikobjektet eller tabellen (markera grafik eller tabell, välj meny Infoga - Bildtext, klicka på OK).  
Därefter går du till stället där referensen ska stå.  
Välj Infoga - Korshänvisning.  
Välj ett av de element för vilka du har definierat en bildtext i listrutan Fälttyp under fliken Referenser.  
Välj t.ex. posten "Illustration" och sedan den illustration som du vill hänvisa till under Urval.  
I listrutan Format väljer du typ av referenspost.  
Till slut klickar du på Infoga.  
Formatet "Över / under" infogar till exempel orden "över "eller "under", oavsett om illustrationen i dokumentet finns ovanför eller nedanför referensen.  
Formatet "Kapitel" förutsätter en kapitelnumrering och en motsvarande formaterad överskrift ovanför illustrationen.  
Formatet "Som sidformatmall" infogar en sidangivelse av den typ som matats in för Numrering under fliken Sida under Format - Sida.  
Referenser har inget stöd i dokument som exporterats till HTML-format.  
Återställa teckenattribut under inmatningen  
När du skriver text och använder direkta formateringar kan du återställa alla formateringar om du vill skriva text i standardformat i stället.  
Skriv texten med de direkta teckenformateringarna, tryck sedan en gång på piltangenten (Högerpil) för att byta tillbaka till standardformatet för stycket.  
Förutsättningen för att detta ska fungera är att du skriver i slutet av det aktuella stycket.  
Exempel  
Du skriver "Detta är", sedan klickar du på ikonerna Fet och Kursiv på textobjektlisten.  
I stället för att klicka på de båda ikonerna igen trycker du en gång på höger piltangent.  
Sedan fortsätter du att skriva i standardformatet för det aktuella stycket.  
Förankra, förstora och förminska fönster  
Ett fönster som Navigator eller Stylist kan du antingen visa som förankrat eller fritt fönster.  
Håll ner Kommando Ctrl -tangenten och dubbelklicka på ett grått område i Navigator-fönstret.  
Navigator-fönstret blir fritt och du kan ställa in storleken genom att dra i kanterna.  
När du är färdig håller du ner Kommando Ctrl -tangenten och dubbelklickar på det gråa området igen, och Navigator förankras vid sin gamla position igen.  
Detsamma gäller för andra förankrade fönster som t.ex. Stylist eller Gallery.  
Söka text med jokertecken  
Öppna dialogrutan Sök och ersätt, t.ex. med Kommando Ctrl +G.  
Markera rutan Reguljärt uttryck.  
Mata in sökordet med eventuella jokertecken och klicka på Sök.  
De reguljära uttrycken anges i en form som bör vara bekant för Unix-användare.  
En stjärna efter ett tecken fungerar som platshållare för ett obestämt antal av tecknet.  
Exempel:  
Om du anger "Hawai*" som sökord så betyder det att ett obestämt antal "i "får, men inte behöver, stå efter "Hawa".  
Orden "Hawa", "Hawai", "Hawaii" hittas.  
En punkt fungerar som platshållare för exakt ett tecken.  
Detta motsvarar jokertecknet? i filnamn.  
För flera tecken som följer direkt efter varandra fungerar kombinationen .* (punkt och stjärna) som platshållare.  
Detta motsvarar jokertecknet * i filnamn.  
Ett styckeslut hittas med dollartecknet ($), det första tecknet i början av ett stycke med kombinationen caret och punkt (^.).  
Det går bara att använda reguljära uttryck inom stycken.  
Det går att använda flera andra jokertecken som finns i en tabellarisk uppställning i %PRODUCTNAME -hjälpen.  
Lista med jokertecken  
Redigera område  
Du kan redigera områdena i ett textdokument genom att välja Format - Områden.  
I den här dialogrutan kan du skydda områden, frige skyddade områden, göra dolda områden synliga, ändra villkor och upphäva områden, d.v.s. omvandla dem till normal text igen.  
Infoga område  
Placera markören på det ställe där du vill infoga ett nytt område, eller markera texten som ska bilda ett område.  
Välj Infoga - Område.  
Du kan göra fler inställningar för området i dialogrutan.  
Klicka på Infoga.  
Då måste rutan Länka markeras.  
I textfältet kan du ange ett filnamn, eller så klickar du på "..." och letar efter en fil i dialogrutan Infoga.  
I kombinationsfältet Område kan du välja ett område i det valda dokumentet.  
När ett dokument öppnas som innehåller länkade områden, tillfrågas du om du vill uppdatera områdena.  
Om du svarar med Ja, så läses de länkade områdena in på nytt.  
Under Windows kan du även använda DDE-mekanismen för att ständigt uppdatera infogade områden så att de har samma status som ursprungsfilerna.  
Områden som filer är möjliga även i HTML-dokument.  
De infogade områdena uppdateras automatiskt när %PRODUCTNAME laddar HTML-dokumentet igen.  
Webbläsare visar områdenas innehåll så som det var när det sparades som HTML-dokument.  
Använda områden  
Områdena i textdokument används till att markera textavsnitt för speciella ändamål.  
Det finns följande områden:  
Områden som textavsnitt med ett annat antal kolumner än den överordnade texten  
Områden som är skyddade för fortsatt redigering  
Områden som bara ska visas när vissa villkor uppfylls eller inte alls  
Områden som ska infogas i ett dokument som filer eller delar av filer  
Områden som när som helst ska överföras till andra textdokument med sin aktuella redigeringsstatus via DDE  
Ett område består alltid av minst ett stycke.  
Om du markerar en text och definierar den som område, avslutas den automatiskt med en styckebrytning.  
Det går även att infoga ett område från ett annat textdokument som område.  
Områden kan också länkas till andra ställen inom ett och samma dokument.  
Om du vill infoga ett nytt stycke direkt före eller efter ett område placerar du markören allra först eller sist i området och trycker på tangenterna Alternativ Alt +Retur.  
Områden och kolumner  
Område med flera kolumner:  
Ett område kan i sin tur innehålla fler områden.  
Denna egenskap gör t.ex. att man kan skapa ett område på en textsida med två kolumner, och definiera ett område med tre kolumner inuti det här området.  
Sida med flera kolumner:  
Sidformateringen, som alltid gäller för alla sidor med den aktualla sidformatmallen, gäller oberoende av områden (Format - Sida - Kolumner).  
Ram med flera kolumner:  
Dessutom kan du infoga ramar, som kan flyttas fritt på sidan, med textkolumner (verktygslist, utrullningslist Infoga, ikon Infoga ram manuellt).  
För de här ramarna kan du t.ex. välja att texten i ramen ska ha ett visst avstånd till ramens kanter (meny Format - Ram, fliken Inramning).  
Även texten utanför ramen kan tilldelas ett avstånd (meny Format - Ram, fliken Textanpassning).  
Språkigenkänning  
Om du har installerat rättstavningen på flera språk så kan %PRODUCTNAME känna igen ord på andra språk och tilldela det rätt språk.  
Förutsättningen är att du inte har markerat rutan Kontrollera alla språk i dialogrutan Verktyg - Alternativ - Språkinställningar - Lingvistik. %PRODUCTNAME kontrollerar i så fall bara i det språk som tilldelats texten som teckenattribut.  
Ord på andra språk framhävs med en röd vågig linje om den automatiska rättstavningskontrollen aktiveras.  
I snabbmenyn till ett sådant ord finns det förslag att det här ordet eller hela stycket ska tilldelas ett av de andra installerade språken, under förutsättning att ordet är rättstavat på respektive språk.  
%PRODUCTNAME kontrollerar rättstavningen för andra språk om du har markerat rutan Kontrollera alla språk i dialogrutan Lingvistik eller om du har tilldelat en text på ett annat språk det riktiga språket som teckenattribut.  
Publicera textdokument som HTML  
%PRODUCTNAME Writer kan, precis som %PRODUCTNAME Calc och %PRODUCTNAME Impress, spara ett strukturerat dokument som webbdokument i HTML-format automatiskt.  
I %PRODUCTNAME Writer väljer du vilka stycken som blir hyperlänkar där dokumentet delas upp i deldokument.  
Grafikobjekt som är inbäddade i dokumentet sparas automatiskt som JPEG-fil i samma katalog som HTML-dokumentet och refereras som IMG-tagg.  
Länkade grafikobjekt bör finnas i samma katalog som HTML-dokumentet så att de kan refereras med en relativ länk.  
Skriv ett textdokument på flera sidor.  
Använd t.ex. mallen Överskrift 2 för överskrifterna till enskilda avsnitt i dokument.  
Välj kommandot Arkiv - Skicka - Skapa HTML-dokument.  
Dialogrutan HTML-dokumentets namn och sökväg öppnas.  
Längst nere i dialogrutan ser du vilken styckeformatmall som fungerar som "avgränsare".  
Om du vill ha en annan styckeformatmall som "avgränsare" väljer du den i kombinationsfältet Akutell formatmall.  
I det här exemplet väljer du Överskrift 2.  
Alla stycken som du har tilldelat den här mallen blir hyperlänkar i HTML-dokumentet.  
Varje hyperlänk öppnar en HTML-sida med underordnat innehåll.  
Ange en sökväg och ett namn för HTML-dokumentet som ska skrivas och klicka på Spara.  
HTML-dokumentet öppnas automatiskt - som alla HTML-dokument skrivskyddat.  
Om du vill redigera det klickar du på ikonen Redigera fil på funktionslisten.  
Så här formaterar du text med kortkommandon medan du skriver  
Så här formaterar du text fet medan du skriver  
Du vill skriva "text i fet stil":  
Skriv "text i" med ett mellanslag efter.  
Tryck på Kommando Ctrl +F.  
Kommando Ctrl +F är kortkommandot för att formatera text fet.  
Skriv "fet".  
Tryck på kortkommandot igen.  
Om du skriver i slutet av ett stycke finns det ett enklare alternativ: tryck en gång på höger piltangent.  
Skriv resten av texten.  
Så här höjer eller sänker du text medan du skriver  
Kortkommandon för textdokument  
Kortkommandon i %PRODUCTNAME  
Dialogruta för rättstavningskontroll  
Dialogrutan öppnas nämligen inte om du väljer Verktyg - Rättstavning - Kontrollera eller trycker på F7 och det inte finns något okänt ord i ditt dokument.  
Då måste du stava ett ord fel eller skriva ett okänt ord med avsikt.  
Dialogrutan Rättstavning visas om du startar rättstavningskontrollen manuellt via menyn eller F7-tangenten.  
Den här metoden har den fördelen att du kan markera en text innan du öppnar dialogrutan och då bara kontrollera stavningen i den här texten.  
Dialogrutan Rättstavning beskrivs utförligt i %PRODUCTNAME -hjälpen.  
Men detta gäller inte om text har markerats, då börjar nämligen kontrollen i början av den markerade texten och slutar där den markerade texten slutar.  
Om rättstavningskontrollen inte börjar i början av dokumentet och når slutet på dokumentet, tillfrågas du i en dialogruta om du vill fortsätta kontrollen i början av dokumentet.  
Först söks alltid de registrerade användarordlistorna igenom.  
Om ordet inte hittas där, söks huvudordlistan igenom.  
Om ordet inte finns där heller, ser du den avbildade dialogrutan där du kan ersätta ordet.  
Skriv det rätt i textfältet eller välj ett i listan med alternativ och klicka sedan på Ersätt.  
Du kan lägga till ordet som står i textfältet Ord i en användarordlista permanent, genom att först välja användarordlistan i kombinationsfältet Ordlista och sedan klicka på kommandoknappen Lägg till.  
Om du har ersatt ordet i textfältet med ett annat kan du kontrollera det andra ordet genom att klicka på Kontrollera ord.  
Om du vill kan du automatiskt lägga till alla okända ord i en text i en aktiverad användarordlista.  
Det finns en beskrivning i %PRODUCTNAME -hjälpen.  
Stänga av punktuppställning eller numrering  
Om %PRODUCTNAME automatiskt fortsätter med en punktuppställning när du trycker på returtangenten trycker du på returtangenten igen om du vill radera punktuppställningstecknet och avsluta punktuppställningen.  
För numreringar gäller motsvarande.  
Om du vill avbryta en numrering som löper över flera stycken med ett stycke utan numrering, raderar du numret framför stycket med Delete-tangenten.  
De följande numren anpassas automatiskt.  
Överföra format i tilldelningsläget  
Så här tilldelar du en ny formatmall i tilldelningsläget:  
Öppna Stylist.  
Markera formatmallen som du vill kopiera i Stylist.  
Klicka på ikonen Tilldelningsläge.  
Peka med musen på objektet som du vill tilldela formatmallen och tryck på musknappen.  
Om du tilldelar en teckenformatmall i tilldelningsläget håller du ner musknappen när du markerar tecknen med musen i stället för att klicka.  
När du vill lämna tilldelningsläget klickar du på ikonen igen eller trycker på Esc.  
Stylist  
Skapa ny formatmall av markering  
Så här skapar du en ny formatmall som kopia av en existerande mall:  
Öppna Stylist.  
Markera en formaterad text eller ett formaterat stycke vars format du vill använda som formatmall.  
Klicka på ikonen i Stylist:  
Ny formatmall av markering  
Du kan också skapa en ny formatmall av markeringen med dra-och-släpp.  
Välj typ av formatmall (styckeformatmallar, teckenformatmallar o.s.v.) genom att klicka på motsvarande ikon överst i Stylist.  
Markera en del av ett stycke eller en text eller ett objekt vars formatering ska ligga till grund för den nya mallen.  
Dra den här delen till huvudområdet i Stylist och släpp musknappen över ett tomt område, d.v.s. när du inte ser någon infogningslinje i Stylist.  
Stylist  
Uppdatera formatmall från markering  
Så här uppdaterar du en formatmall:  
Öppna Stylist.  
I dokumentet markerar du en formaterad text eller ett formaterat stycke vars format du vill använda som formatmall.  
I Stylist markerar du formatmallen som ska uppdateras (klicka enkelt, dubbelklicka inte!)  
Klicka på ikonen i Stylist:  
Uppdatera formatmall  
Du kan också uppdatera formatmallen med dra-och-släpp.  
I Stylist markerar du mallen som du vill uppdatera.  
Markera en del av texten i stycket vars format du nu vill använda till mallen som är markerad i Stylist.  
Dra textdelen till huvudområdet i Stylist och släpp musknappen över en post, d.v.s. när du ser infogningslinjen i Stylist.  
Styckeformatmallen som står direkt ovanför infogningslinjen får det nya formatet.  
Stylist  
Upphöjd och nedsänkt text  
Det finns följande möjligheter att höja och sänka text:  
Använd kortkommandona Ctrl+H och Ctrl+T.  
Använd kommandot Format - Tecken - Position.  
Använd ikonerna: öppna snabbmenyn på textobjektlisten, välj Synliga knappar och markera Nedsänkt och Upphöjt på undermenyn.  
Nu visas ikonerna på textobjektlisten.  
Så här höjer eller sänker du text medan du skriver  
Du vill skriva 1 m² med upphöjd tvåa:  
Skriv 1 m2.  
Efter 2 trycker du på mellanslagstangenten eller en annan tangent som definierar ett ordslut.  
Av m2 blir det automatiskt m² om det här ersättningsparet finns under fliken Ersättning under Verktyg - AutoKorrigering / AutoFormat.  
Du kan utvidga listan så mycket du vill.  
Fortsätt att skriva normalt efter den automatiska ersättningen.  
Du vill skriva H2O med nedsänkt tvåa:  
Skriv H:et.  
Tryck på Kommando Ctrl +T.  
Kommando Ctrl +T är kortkommandot för nedsänkt text, Kommando Ctrl +H för upphöjd text.  
Skriv 2.  
Tryck på kortkommandot igen.  
Om du skriver i slutet av ett stycke finns det ett enklare alternativ: tryck en gång på höger piltangent.  
Skriv O.  
Formatera text upphöjd eller nedsänkt i efterhand  
Du vill t.ex. omvandla texten H2O till H2O med nedsänkt tvåa i efterhand.  
Använd tangentkombinationen som beskrivs ovan eller gör på följande sätt:  
Markera tecknet som du vill höja eller sänka.  
I det här exemplet markerar du 2:an.  
Välj Format - Tecken.  
Dialogrutan Tecken öppnas.  
Klicka på fliken Position.  
Välj alternativet Nedsänkt och klicka på OK.  
2:an är nu nedsänkt.  
Format - Tecken - Position  
Verktyg - AutoKorrigering / AutoFormat - Ersättning  
Infoga eller radera rader / kolumner via tangentbordet  
Om du vill infoga eller radera rader och kolumner via tangentbordet gör du så här:  
Om du vill infoga en ny kolumn eller rad växlar du först till infogningsläget för tabeller med tangentkombinationen Alternativ Alt +Insert.  
Detta gäller i tre sekunder, och under den tiden kan du trycka på respektive piltangent för att infoga en ny rad eller kolumn till höger, vänster, ovanför eller nedanför den aktuella raden eller kolumnen.  
Om du dessutom håller ner Kommando Ctrl -tangenten samtidigt som piltangenten, så delas den intilliggande cellen.  
Om du vill radera en kolumn eller rad växlar du först till raderingsläget för tabeller med tangentkombinationen Alternativ Alt +Delete.  
Detta gäller i tre sekunder, och under den tiden kan du trycka på respektive piltangent för att radera en rad eller kolumn till höger, vänster, ovanför eller nedanför den aktuella raden eller kolumnen.  
Om du håller ner Kommando Ctrl -tangenten samtidigt som piltangenten, så sammanfogas den aktuella cellen med den intilliggande cellen till en cell.  
Radera tabell  
Om du vill radera en hel tabell i ett textdokument har du följande möjligheter:  
Markera från slutet av stycket före tabellen till början av stycket efter tabellen.  
Tryck på Delete-tangenten eller backstegstangenten.  
Eller sätt markören i tabellen, markera alla celler, t.ex. med Kommando Ctrl +A, öppna snabbmenyn och välj Rad - Radera.  
Den här metoden går också att använda i början eller slutet av dokumentet.  
Infoga tabell  
Det finns olika sätt att infoga en tabell i ett textdokument:  
Infoga en tom tabell med musen  
Placera markören på det ställe i texten där du vill infoga tabellen.  
Peka med musen på ikonen Infoga tabell på utrullningslisten Infoga.  
Tryck på musknappen och dra musen nedåt och åt höger tills du har markerat så många rader och kolumner som du behöver i förhandsvisningsfältet.  
Släpp sedan musknappen. (Om du vill avbryta processen drar du musen uppåt eller åt vänster innan du släpper musknappen tills du ser att det står Avbryt i förhandsvisningsfältet.)  
Infoga en tom tabell via dialogruta  
Placera markören på det ställe i texten där du vill infoga tabellen.  
Klicka kort på ikonen Infoga tabell på utrullningslisten Infoga.  
Dialogrutan Infoga tabell visas.  
Infoga från %PRODUCTNAME Calc via urklippet  
Öppna ditt textdokument och ett %PRODUCTNAME Calc-dokument som innehåller ett cellområde som du vill klistra in i textdokumentet.  
Markera ett cellområde i tabelldokumentet.  
Kopiera det till urklippet, t.ex. med Ctrl+C.  
Byt till textdokumentet.  
Nu har du olika möjligheter att klistra in cellområdet:  
Om du väljer det "normala" kommandot Redigera - Klistra in eller Ctrl+V klistrar du in cellområdet som OLE-objekt.  
Du kan dubbelklicka på OLE-objektet och sedan redigera det med verktygen och kommandona från %PRODUCTNAME Calc.  
Klicka utanför objektet när du vill lämna redigeringsläget.  
Om du väljer Redigera - Klistra in innehåll öppnas dialogrutan Klistra in innehåll där du väljer bland flera möjligheter.  
Samma möjligheter finns också på undermenyn till ikonen Klistra in på funktionslisten:  
Urval  
Klistras in som...  
"%PRODUCTNAME 6.0-tabell" resp. "Star Embed Source "  
OLE-objekt - som med Ctrl+V eller dra-och-släpp  
GDI-metafil  
Grafik  
Bitmap  
Grafik  
HTML  
HTML-tabell  
Oformaterad text  
Bara text, tabbar som avgränsare  
Formaterad text [RTF]  
Texttabell  
DDE-länk (bara i Windows)  
Tabellstruktur och innehåll, utan formatering.  
Med uppdatering  
Klistra in från %PRODUCTNAME Calc med dra-och-släpp  
Öppna ditt textdokument och ett %PRODUCTNAME Calc-dokument som innehåller ett cellområde som du vill klistra in i textdokumentet.  
Markera ett cellområde i tabelldokumentet.  
Klicka på det markerade cellområdet och håll ner musknappen.  
Fortsätt att hålla ner musknappen och vänta ett ögonblick.  
Dra det markerade cellområdet till textdokumentet utan att släppa musknappen.  
Om textdokumentet inte är synligt måste du först föra muspekaren till textdokumentets symbol på aktivitetsfältet och vänta ett ögonblick tills textdokumentet öppnas.  
I textdokumentet följer en grå infogningsmarkör muspekaren och visar var tabellen kan placeras.  
Släpp musknappen när den gråa infogningsmarkören visar var tabellen ska klistras in.  
Anpassa tabellbredd  
Tabellens beteende påverkas av tabellens förinställning, som du gör i dialogrutan Verktyg - Alternativ - Textdokument - Tabell eller genom att klicka på motsvarande ikoner på tabellobjektlisten.  
Du kan här välja mellan fast, fast / proportionell och variabel.  
Tabelläge fast innebär att när man gör en cell bredare blir den intilliggande cellen i motsvarande mån smalare.  
Andra celler påverkas inte, tabellbredden förblir densamma.  
Tabelläge fast och proportionell innebär att samtliga intilliggande celler i motsvarande riktning förminskas, breda celler proportionellt mer än smala.  
Tabellbredden förblir densamma.  
Tabelläge variabel innebär att hela tabellens bredd är variabel - hela tabellen blir helt enkelt bredare när en cell görs bredare.  
Även vid infogning och radering avgör tabelläget hur intilliggande celler, rader eller kolumner ska påverkas.  
I fast läge infogas bara nya rader och kolumner om det finns plats.  
Upprepa flera överskriftsrader i tabeller  
Om du vill att mer än en rad ska upprepas automatiskt i en tabell vid sidbrytning gör du så här:  
Markera hela den första raden i tabellen.  
Öppna snabbmenyn och välj Cell - Dela.  
I dialogrutan Dela celler väljer du "horisontellt" som riktning.  
Ange antalet rader som ska upprepas och bekräfta med "OK".  
Efter en sidbrytning upprepas nu alla rader som har skapats på det här sättet i början av tabellen.  
Förstora och förminska celler i en texttabell  
Du kan ändra bredden och höjden på rader och kolumner via tangentbordet, genom att dra med musen eller genom att använda kommandon på snabbmenyn.  
Kolumnbredden kan också ändras numeriskt via en dialogruta.  
Du uppnår dessutom en jämn fördelning med ikonerna på utrullningslisten Optimera på tabellobjektlisten.  
Med hjälp av musen kan du ändra raderna och kolumnerna i tabellen eller på linjalerna.  
Peka på en skiljelinje i tabellen, så blir muspekaren till en skiljesymbol.  
Håll nu ner musknappen och dra så flyttas linjen. (Eventuellt måste du klicka en gång utanför tabellen innan den här metoden fungerar.) På samma sätt kan du flytta de skiljelinjer som är synliga på linjalerna.  
När du förstorar och förminskar med hjälp av tangentbordet måste du alltid hålla ner Alternativ Alt -tangenten.  
Hur mycket kan du ställa in separat för rader och kolumner i dialogrutan Verktyg - Alternativ - Textdokument - Tabell i området Tangentbordshantering.  
Den aktuella raden eller kolumnen förstoras eller förminskas i högra eller nedre kanten.  
Tryck på Alternativ Alt -tangenten och skifttangenten samtidigt, så flyttas den vänstra eller övre kanten.  
Två exempel:  
Sätt markören mitt i en större texttabell.  
Håll ner Alternativ Alt -tangenten och tryck på den högra piltangenten.  
Den aktuella kolumnen blir så mycket bredare som är inställt vid Flytta / Kolumn under Verktyg - Alternativ... - Textdokument - Tabell.  
Kolumnens vänstra kant stannar kvar på sin plats, högra kanten flyttas.  
Håll ner Alternativ Alt -tangenten tillsammans med skifttangenten och tryck på den högra piltangenten.  
Nu stannar högra kanten kvar på sin plats och vänstra kanten flyttas åt höger.  
Kolumnen förminskas alltså.  
För riktningen uppåt / nedåt gäller motsvarande, men raderna är enligt förinställningen redan minimalt höga, vilket innebär att du först måste förstora dem innan du kan se en effekt som liknar den hos kolumnerna.  
Om du dessutom håller ner Kommando Ctrl -tangenten, gäller förstoringen eller förminskningen bara för den aktuella cellen istället för hela raden eller kolumnen.  
Måtten för hela tabellen förblir nu fasta.  
Skapa dokumentmall  
För att dina användardefinierade stycke - eller teckenformatmallar ska vara tillgängliga även i andra dokument skapar du en dokumentmall.  
Dokumentmallen innehåller alla formatmallar som finns i det aktuella dokumentet.  
Om du vill kan du radera alla texter från det aktuella dokumentet så att bara mallarna finns kvar.  
Du kan använda formatmallarna från ett textdokument i ett annat textdokument: meny Format - Mallar - Ladda.  
Välj Arkiv - Dokumentmall - Spara.  
I dialogrutan Dokumentmall väljer du kategorin där dokumentmallen skall sparas.  
I textfältet Ny dokumentmall anger du namnet på dokumentmallen.  
Klicka på OK.  
Senare kan du öppna en dialogruta under Arkiv - Nytt - Mallar och dokument där du kan välja ut din dokumentmall.  
Ett nytt dokument öppnas som är en kopia av dokumentmallen.  
Dina stycke - och teckenformatmallar är tillgängliga i det nya dokumentet.  
Arkiv - Dokumentmall - Spara  
Definiera standardmall  
Om du märker att du måste ändra formateringarna i dina nya dokument varje gång för att anpassa utseendet på sidorna efter dina önskemål kan du använda en egen mall, den så kallade Standardmallen.  
Den här standardmallen används alltid om du öppnar ett nytt textdokument, t.ex. via Arkiv - Nytt - Textdokument.  
Skapa eller öppna ett dokument som innehåller alla formatmallar med de formateringar som du föredrar.  
Om du vill kan du radera innehållet i dokumentet så att bara formatmallarna och andra inställningar finns kvar.  
Spara dokumentet som mall med Arkiv - Dokumentmall - Spara i kategorin Standard.  
Då sparas dokumentet som mall i katalogen {installpath} / user / template {installpath }\user\template.  
Välj Arkiv - Dokumentmall - Administrera.  
Dubbelklicka på "Standard" i den vänstra listrutan där dokumentmallarna är listade.  
Under posten "Standard" ser du nu namnet på malldokumentet som du har sparat.  
Klicka på den.  
Välj Definiera som standardmall på snabbmenyn.  
Stäng dialogrutan.  
Nu används malldokumentet som ny standardmall.  
Återställa standardmall  
Välj Arkiv - Dokumentmall - Administrera.  
Öppna snabbmenyn i en av listrutorna eller öppna undermenyn till kommandoknappen Kommandon.  
Välj Återställ standardmall.  
Då öppnas en undermeny där alla dokumenttyper finns angivna för vilken du har valt en egen standardmall.  
Välj den dokumenttyp som du vill tilldela den förinställda standardmallen igen.  
Dokumentmallar och formatmallar  
Dokumentmallarna i %PRODUCTNAME är filer som du kan använda som utgångspunkt för dina egna dokument.  
Dokumentmallarna kan innehålla texter, logotyper, andra grafiska objekt med mera.  
Dessutom innehåller varje dokumentmall ett flertal formatmallar som du kan titta på i Stylist.  
Standardmallen används alltid när du skapar ett nytt (oftast tomt) dokument via t.ex. Arkiv - Nytt.  
Det finns malltyper för nästan alla dokumenttyper.  
I %PRODUCTNAME -hjälpen till textdokument finns det en lista med de olika mallarna för textdokument, motsvarande gäller för mallarna till presentationsdokument och tabelldokument.  
Om du väljer Format - Mallar - Katalog visas en dialogruta som innehåller olika formatmallar för redigering beroende på av vilken typ det aktuella dokumentet är.  
Om du t.ex. har öppnat ett textdokument och väljer det här kommandot, ser dialogrutan ut så här:  
Här kan du, ungefär som i Stylist, välja typ av formatmall i en listruta, ändra mallarna som hör till den här typen, radera mallar som du själv har skapat och skapa nya mallar.  
Men du kan också klicka på Administrera.  
Då visas en dialogruta med ett innehåll som liknar innehållet på följande bild:  
I den här dialogrutan kan du kopiera formatmallarna, som finns i en viss dokumentmall eller i ett visst dokument, en och en till ett annat dokument.  
Titta på bilden.  
Om du dubbelklickar på ett mappnamn i det vänstra fönstret visas alla dokumentmallar som finns i mappen.  
Om du dubbelklickar på en sådan fil ser du de båda områdena Mallar och Konfiguration.  
Även här kan du öppna respektive lista med objekt genom att dubbelklicka.  
Men för ett dokument ser du bara mallarna som verkligen används i respektive dokument.  
Om du drar element från en dialogsida till en annan med dra-och-släpp, ser du hur muspekaren signalerar var du kan placera innehållet.  
Antingen är muspekaren en genomstruken cirkel - då kan du inte placera innehållet på muspekarens plats - eller så har muspekaren en infogningslinje som anger platsen där innehållet placeras när du släpper musknappen.  
Justera text längs linje  
Justera text längs frihandslinje  
Rita frihandslinjen (utrullningslist Ritfunktioner).  
Dubbelklicka på linjen.  
Skriv den önskade texten eller kopiera den från urklippet.  
Välj Format - FontWork.  
Klicka t.ex. på ikonen Rotera.  
Justera text längs rät linje  
Om du vill snedställa en text så att den löper exakt från en punkt på textsidan till en annan, gör du så här:  
Rita en rät linje från den ena punkten till den andra med hjälp av ritfunktionerna.  
Välj linjenstilen "Osynlig" i listrutan på objektlisten.  
Dubbelklicka på den nu osynliga linjen (de båda punkterna i varje ände syns fortfarande: dubbelklicka precis mittemellan dem).  
Mata in texten och klicka sedan utanför linjeobjektet.  
Använda animerad text  
Gör så här:  
1.  
Öppna ett nytt tomt %PRODUCTNAME Writer-dokument.  
2.  
Välj en bakgrund för hela sidan under Format - Sida.  
3.  
Öppna utrullningslisten Ritfunktioner på verktygslisten och klicka på ikonen Rektangel.  
4.  
Rita upp en rektangel mitt på sidan:  
5.  
Öppna snabbmenyn till det markerade ritobjektet.  
6.  
Välj Yta för att ge rektangelns yta en annan färg.  
7.  
Välj alternativet Färggradient till vänster under fliken Yta och välj till exempel "Färggradient 4".  
Stäng dialogrutan med OK.  
8.  
Öppna snabbmenyn igen och välj Linje....  
Här kan du bestämma egenskaperna för rektangelns inramning.  
9.  
Välj en färg och bredd för linjen.  
Stäng dialogrutan med OK.  
10.  
Dubbelklicka i mitten av rektangeln.  
Nu kan du skriva in en text.  
Det gör ingenting om texten är bredare än rektangeln.  
11.  
Öppna sedan snabbmenyn och välj Text.  
12.  
I dialogrutan Text klickar du på fliken Animerad text.  
Välj alternativet "Genomlöpa" i kombinationsfältet i området Effekter animerad text.  
Under fliken Text kan du ställa in avståndet från ramen till vänster och höger. (Ramens kant går till hälften inåt och till hälften utåt.) Klicka på OK.  
13.  
Nu behöver du bara avmarkera rektangeln genom att klicka på ett annat ställe i dokumentet.  
Texten börjar genast att rulla.  
14.  
Om du vill ändra storleken på den animerade texten, markerar du rektangeln igen och dubbelklickar i mitten.  
Nu kan du markera texten och till exempel tilldela den en större teckenstorlek.  
Du kan förstora vyn genom att antingen välja Visa - Skala... eller genom att öppna snabbmenyn till fältet som visar skalan i statuslisten (eller dubbelklicka i fältet).  
Om bildskärmsvisningen skall uppdateras använder du tangentkombinationen Skift + Kommando Ctrl +R.  
Skriva text med stora eller små bokstäver  
Hur kan text formateras om till bara stora eller små bokstäver?  
Du har följande möjligheter att formatera om text till stora eller små bokstäver.  
Bestäm om texten bara ska få en teckeneffekt för visning och utskrift eller om tecknen ska ersättas permanent:  
Stora bokstäver: markera text, välj Format - Tecken, klicka på fliken Teckeneffekt och välj effekten Versaler.  
Små bokstäver: markera text, välj Format / Tecken, klicka på fliken Teckeneffekt och välj effekten Gemener.  
Omvandla till stora bokstäver: markera text, välj Format - Bokstäver / tecken - Stora bokstäver.  
Omvandla till små bokstäver: markera text, välj Format - Bokstäver / tecken - Små bokstäver.  
Centrera text vertikalt på sidan  
Om du vill centrera en text vertikalt mellan övre och undre sidmarginalen gör du så här:  
1.  
Markera texten.  
2.  
Klicka på ikonen Infoga ram manuellt på utrullningslisten Infoga uppe på verktygslisten.  
3.  
Rita upp en ram på sidan.  
Den markerade texten sätts automatiskt i ramen.  
4.  
Formatera texten och dimensionera ramens storlek så att den omger texten så tätt intill som möjligt.  
Om du vill formatera texten måste du först markera den.  
Upphäv markeringen av ramen genom att klicka en gång utanför ramen och sedan direkt i texten.  
När du vill markera själva ramen igen klickar du på ramens kant.  
5.  
Öppna ramens snabbmeny och ändra föränkringen till "Vid sidan".  
6.  
Du kan nu dra textramen med musen vart du vill på sidan.  
Du kan också använda ikonerna i objektlisten för att placera ramen horisontellt och / eller vertikalt vid en marginal eller i mitten.  
7.  
I dialogrutan kan du redigera den markerade ramens egenskaper.  
8.  
Ta bort ramens kant under fliken Inramning i dialogrutan Ram, annars skrivs den ut tillsammans med dokumentet.  
Klicka på symbolen helt utan linjer längst till vänster i området Linjeplacering.  
Då har ramen inte kvar kanten som kan skrivas ut.  
Om du vill välja bort den gråa kanten som du kan se på bildskärmen, men som inte skrivs ut, använder du menykommandot Visa - Textbegränsningar.  
Inmatning av text på valfritt ställe  
Med direktmarkören kan du skriva in text var som helst på sidan i ditt textdokument.  
1.  
Klicka på ikonen (Direktmarkör på / av) på verktygslisten.  
Med den här ikonen sätter du på och stänger av direktmarkören.  
Om ikonen är intryckt visar det att direktmarkören aktiverad.  
2.  
Klicka på ett tomt ställe i textdokumentet.  
Muspekarens form visar hur den inmatade texten justeras.  
Vänsterjusterat  
Centrerat  
Högerjusterat  
3.  
Mata in den önskade texten. %PRODUCTNAME sätter automatiskt in det antal tomma rader, tabbar och mellanrum som behövs.  
Infoga externt textdokument  
Om du vill infoga text från ett annat textdokument i det aktuella textdokumentet, finns det flera olika möjligheter:  
Du kan kopiera den externa texten till urklippet och klistra in den i det aktuella dokumentet.  
Detta är snabbt och enkelt men om det externa dokumentet ändras i efterhand visas inte det i det aktuella dokumentet.  
Du kan infoga den externa texten som länk.  
Den externa texten infogas som länk i området.  
Fördelen är att ändringar i det externa dokumentet nästan automatiskt visas i det aktuella dokumentet.  
Om du infogar den externa texten i en textram har du redan innan den externa texten är färdig kontrollen över placeringen av texten på din sida - vilket t.ex. är viktigt om du gör en egen tidning.  
Med länkade ramar kan du bestämma hur den externa texten ska fördelas över flera sidor.  
Om du vill ha texten i ramar ritar du upp ramarna med musen (verktygslisten, utrullningslisten Infoga, ikonen Ram).  
Om du vill ha texten i flera länkade ramar, så ritar du upp alla dessa ramar.  
Om du arbetar med länkade ramar där texten automatiskt löper från en ram till nästa, så definierar du nu länkningen (ikonen Länka på objektlisten).  
Placera textmarkören på det ställe där den externa texten ska börja.  
Välj Infoga - Område....  
Dialogrutan Infoga område visas.  
Markera fältet Länk.  
Nu kan du klicka på Välj ut och välja det externa textdokumentet.  
Om det innehåller namngivna områden, så kan du välja ut ett av dem i kombinationsfältet Område, i annat fall infogas hela dokumentet.  
Mata in ett eget namn för området i textfältet.  
Det här namnet visas t.ex. i Navigator.  
Klicka på Infoga och stäng dialogrutan med stängningsknappen.  
Det externa textdokumentet har infogats som länkat område.  
Förbinda textdokument  
Så bifogar du ett dokument till ett textdokument.  
Placera markören i slutet av det första dokumentet och välj meny Infoga / Fil....  
Välj ut dokumentet som skall laddas i dialogrutan och ladda det.  
Dokumentet infogas nu i slutet av det första dokumentet.  
Framhäva text  
Du har många olika möjligheter att framhäva text.  
Här nämner vi några:  
Utforma texten i fetstil eller i ett annat teckensnitt, ändra textens färg och bakgrund, centrera texten, bara för att nämna några av möjligheterna.  
Om du vill framhäva ett helt stycke optiskt, öppnar du snabbmenyn och väljer Stycke och t.ex. fliken Inramning.  
Här kan du välja ut en inramning som ramar in stycket, med skugga om du vill det.  
Ändra eventuellt avstånden mellan inramning och stycketext i området Avstånd till innehåll.  
Du kan länka samman textramarna om texten skall löpa vidare från en ram till nästa.  
Tilldela stycket en bakgrundsfärg (via Format - Stycke - Bakgrund).  
Använd ritfunktionen Text: med ikonen Text på utrullningslisten Ritfunktioner (till vänster på verktygslisten) ritar du upp en ram och infogar text.  
Den här texten kan du placera var du vill, rotera den i valfria vinklar eller placera den i kurvor med Format - FontWork och tippa bokstäverna.  
Format - FontWork  
Mata in ny text  
Så här matar du in ny text:  
Öppna ett textdokument eller skapa ett nytt.  
Mata in text via tangentbordet.  
Om du vill använda specialtecken som inte finns på ditt tangentbord väljer du Specialtecken på menyn Infoga och väljer tecken i dialogrutan.  
Tryck på returtangenten när du ska börja ett nytt stycke.  
Radslut  
Du behöver inte bekymra dig om radsluten eftersom programmet automatiskt styr radbrytningen.  
Du trycker bara på returtangenten när du vill inleda ett nytt stycke.  
Korrigera automatiskt  
Det innebär t.ex. att alla meningar automatiskt börjar med stor bokstav.  
Komplettera ord  
Du har också hjälp av den automatiska kompletteringen av ord när du skriver:  
Om du skriver in ett längre ord upprepade gånger, föreslår %PRODUCTNAME Writer det här ordet.  
Tryck på returtangenten för att acceptera förslaget.  
Ordkomplettering  
Infoga, redigera och länka textramar  
Infoga textram  
Sätt texten i en textram.  
Om du vill föra över text till en textram gör du på följande sätt:  
1.  
Markera texten som ska vara i ramen.  
2.  
Den heter Infoga ram manuellt.  
Släpp musknappen direkt på ikonen eller klicka kort på ikonen när du ser utrullningslisten som fönster.  
Om du håller ner musknappen och drar neråt från ikonen kan du fortsätta att hålla ner musknappen och välja ett antal kolumner.  
Släpp musknappen när du har valt ut önskat antal kolumner.  
3.  
När du nu flyttar muspekaren i textdokumentet har den ändrat sin form till ett hårkors.  
Det visar att du nu kan rita upp en ram.  
Om du inte vill göra det trycker du på Esc-tangenten för att förvandla muspekaren till en markör igen.  
4.  
Använd hårkorset för att rita upp en ram som visar den nya platsen för stycket.  
Den markerade texten klipps nu automatiskt ut från den normala texten och klistras in i textramen.  
Du kan klicka på textramens kant om du vill markera den.  
En markerad textram känner du igen på de åtta handtagen, fyra i hörnen och en i mitten av varje ramlinje.  
Redigera textram  
Om en textram är markerad, kan du förändra den genom att hålla ner musknappen och dra.  
Om du drar i kanten utanför ett handtag så flyttas hela ramen.  
Om du drar i ett av handtagen, ändras ramens storlek.  
Det motsatta hörnet eller den motsatta sidan till handtaget stannar kvar på sin plats.  
Genom att dra i ett handtag på en sida sträcker eller krymper du textramen i bara en riktning, medan du kan förstora eller förminska den i båda dimensioner genom att dra i ett handtag i ett hörn.  
Om du håller ner skifttangenten när du drar i ett av de åtta handtagen, ändras ramens storlek proportionellt, alltså med samma sidförhållande.  
Du kan göra fler inställningar genom att öppna snabbmenyn till den aktiverade textramen.  
På snabbmenyn till en textram kan du till exempel välja Justering i förhållande till andra ramar, ritobjekt och grafik med mera.  
Med undermenyn Textanpassning väljer du om och på vilken sida av textramen den normala löpande texten finns i ditt dokument.  
Om du klickar på Ram på snabbmenyn, motsvarar det menykommandot Format - Ram.  
Det öppnar en dialogruta som gör alla egenskaper för ramen tillgängliga.  
I textramen står samma funktioner till förfogande som vid textdokument: textramar kan till exempel förutom texten även innehålla grafik, ha flera kolumner och så vidare.  
Länka textramar  
Du kan koppla ihop flera textramar med varandra, även på olika sidor i dokumentet.  
Då löper texten automatiskt från en ram till nästa.  
1.  
Om du vill länka ihop ramar, klickar du på kanten på den ram som du vill länka ihop med en annan ram.  
Åtta handtag visas på kanten.  
2.  
Klicka på ikonen Länka på objektlisten.  
3.  
Klicka på ramen som ska länkas.  
Om en länkad ram är markerad visas länkningarna med en linje på bildskärmen.  
När en ram länkas ihop med en efterföljande ram så fixeras höjden automatiskt.  
Höjden anpassas sedan inte mer till ramens innehåll automatiskt.  
Det är bara den sista ramen i en kedja som kan anpassa sin höjd till textinnehållet.  
När du har markerat en ram och klickar på ikonen Länka på objektlisten, ändras muspekarens utseende.  
Den kan nu visa två symboler: en kedja med pil om det är möjligt att länka ihop två ramar med musen, eller en kedja med stoppskylt om det inte är möjligt att länka ihop ramar vid den aktuella positionen.  
I statuslisten visas alltid en informationstext, t.ex. varför det inte är möjligt att länka.  
Det är bara möjligt att göra en länkning från en ram till nästa.  
Det betyder att en ram som redan är länkad till en annan ram inte kan länkas ihop med ytterligare en ram.  
Därför kan ikonen "Länkning" inte aktiveras om en ram redan har en följande ram.  
Dessutom är det bara möjligt att öppna länkningen av två ramar från den föregående ramens håll med ikonen Lös upp länkning.  
Att länka ihop ramar är inte tillåtet om följande villkor är uppfyllda:  
Målet är inte tomt.  
En (automatiskt) etiketterad ram är inte tom och kan därför inte vara mål för en länkning.  
Målet har redan en föregående ram.  
Källa och mål står i olika områden, t.ex. en ram i ett sidhuvud och en ram i en sidfot.  
Källan har redan en följande ram.  
Källa och mål är identiska.  
Slutna kedjor eller kedjor inifrån och utåt eller utifrån och inåt är inte heller tillåtna.  
Ett exempel på det sistnämnda är om du har infogat en ram i en annan och vill länka ihop dem med varandra.  
Infoga text  
Öppna ett dokument som redan finns.  
Placera markören med hjälp av musen eller med piltangenterna på det ställe där texten ska läggas till och mata sedan in ny text.  
Textdokumentet är som regel i infogningsläge; texten som kommer efter infogningsstället flyttas framåt när du skriver den nya texten.  
Om du vill att texten som kommer efter infogningsstället ska skrivas över av den nya texten väljer du överskrivningsläget.  
Navigera och markera med tangentbordet  
Använd piltangenterna och tangenterna Home, End, Page Up och Page Down när du navigerar och markerar med tangentbordet.  
Några tangenter har olika funktioner beroende på om bara de används eller om de används tillsammans med Kommandotangenten Ctrl-tangenten.  
Följande tabell är en översikt över tangenternas funktioner för navigering.  
Tangent  
Funktion  
+ Kommandotangent Ctrl-tangent  
Piltangenter höger / vänster  
gå ett tecken åt vänster eller höger  
ett ord åt vänster eller höger  
Piltangenter upp / ned  
gå en rad uppåt eller nedåt  
flytta det aktuella stycket uppåt eller nedåt  
Home  
gå till början av den aktuella raden  
gå till början av dokumentet  
Home  
i en tabell  
gå till början av den aktuella cellen  
1. gå till början av den aktuella cellen  
2. gå till början av tabellen  
3. gå till början av dokumentet  
End  
gå till slutet av den aktuella raden  
gå till slutet av dokumentet  
End  
i en tabell  
gå till slutet av den aktuella cellen  
1. gå till slutet av den aktuella cellen  
2. gå till slutet av tabellen  
3. gå till slutet av dokumentet  
Page Up  
bläddra en bildskärmssida uppåt  
byta till sidhuvudet och tillbaka  
Page Down  
bläddra en bildskärmssida nedåt  
byta till sidfoten och tillbaka  
Rotera text  
Om du vill rotera text matar du in den i en textteckenram:  
Öppna utrullningslisten Ritfunktioner på verktygslisten.  
Klicka på ikonen Text på utrullningslisten.  
Muspekaren visar att du kan rita upp en textteckenram.  
Rita upp en textteckenram, släpp musknappen och mata in texten.  
Klicka på kanten av textteckenramen.  
Teckenobjektlisten visas på vilken ikonen Objekt-rotationsläge finns.  
Klicka på ikonen.  
Om du nu klickar på ett av handtagen i hörnorna på textteckenramen och drar musen roteras hela ramen med texten.  
På snabbmenyn till textramen kan du öppna dialogrutan Position och storlek där fliken Rotation finns.  
Här kan du definiera rotationsvinkeln.  
Ritfunktioner - Text  
Markera och radera text  
Radera ett tecken  
Om markören står efter tecknet som ska raderas, trycker du på backstegstangenten (ovanför returtangenten).  
Den här tangenten raderar ett tecken till vänster om markören.  
Om markören står framför tecknet som ska raderas trycker du på Delete-tangenten (ovanför piltangenterna).  
Den här tangenten raderar ett tecken till höger om markören.  
Radera texter  
Markera texten som ska raderas med musen  
Klicka med vänster musknapp på det första tecknet som ska raderas.  
Håll ner musknappen och dra till det sista tecknet som ska raderas.  
Släpp musknappen.  
Tryck på Delete-tangenten för att radera den markerade texten.  
Markera texten som ska raderas med tangentbordet  
Placera markören framför det första tecknet som ska raderas.  
Tryck på skifttangenten.  
Flytta markören med hjälp piltangenterna och placera den efter det sista tecknet som ska raderas.  
Släpp skifttangenten.  
Texten markeras.  
Tryck på Delete-tangenten för att radera den markerade texten.  
Om du inte raderar texten med Delete-tangenten utan med tangentkombinationen Kommando Ctrl +X, klipps texten ut och placeras i urklippet.  
Du kan då klistra in den på andra ställen igen, t.ex. med tangentkombinationen Kommando Ctrl +V.  
Radera texter som inte hänger ihop  
Tryck på Kommando Ctrl -tangenten och håll ner den.  
Klicka med den vänstra musknappen på det första tecknet i den första texten som ska raderas.  
Håll ner musknappen och dra till det sista tecknet i den här texten.  
Släpp musknappen och Kommando Ctrl -tangenten.  
Upprepa steg 1 till 4 för varje text som ska raderas.  
Tryck på Delete-tangenten för att radera de markerade texterna.  
Fotnoter och slutnoter  
I ditt textdokument kan du visa fotnoter i slutet av sidan (eller av kolumnen vid layout med flera kolumner) eller i slutet av dokumentet.  
Inställningarna väljer du med Verktyg - Fotnoter.  
Följande information gäller även för slutnoter.  
Slutnoter är fotnoter som samlas i slutet av ett dokument i stället för längst ned på sidan.  
Du kan enkelt hoppa från ett fotnotsankare i dokumentet till fotnotstexten genom att klicka på fotnotsankaret.  
Med tangenten PageUp kommer du tillbaka till texten från fotnoten.  
Du kan påverka fotnoternas format genom att ändra styckeformatmallen "Fotnot", som automatiskt används för fotnoterna.  
Om du vill radera en fotnot räcker det att radera fotnotsmärket i texten.  
Fotnotstexten raderas då automatiskt.  
Avstavning  
Du kan göra avstavningen i textdokument automatiskt eller manuellt.  
Den automatiska avstavningen är ett attribut i stycken och styckeformatmallar.  
Det betyder att du kan sätta på eller stänga av avstavningen för ett stycke eller för ett styckeformat och välja egenskaper för avstavningen.  
Den manuella avstavningen gör det möjligt att styra individuellt hur ord avstavas, men tar därför också mycket tid.  
Den automatiska avstavningen  
Standardinställningen är att den automatiska avstavningen är aktiverad.  
Om du vill aktivera avstavningen för ett eller flera markerade stycken, öppnar du snabbmenyn och väljer Stycke.  
Om du vill aktivera avstavningen för alla stycken som är formaterade med en viss styckeformatmall, öppnar du snabbmenyn på ett sådant stycke och väljer Redigera styckeformatmall.  
Om du vill använda avstavningen för alla stycken redigerar du styckeformatmallen Standard som de andra styckeformatmallarna bygger på.  
I dialogrutan som öppnas klickar du på fliken Textflöde.  
I området Avstavning markerar du rutan Automatisk.  
Den manuella avstavningen  
Om du vill göra en manuell avstavning, placerar du textmarkören på det ställe i ordet där det ska avstavas och trycker på Kommando Ctrl -.  
Ordet avstavas om det är möjligt, även om den automatiska avstavningen är avstängd för stycket.  
Om du har matat in en avstavning manuellt använder %PRODUCTNAME inte de följande automatiska avstavningarna i det här ordet.  
An-tarcti-ca.  
Du vill nu avstava ordet på följande sätt:  
Ant-arc-ti-ca.  
Du matar in alla tre avstavningarna manuellt, även den sista framför "ca".  
Det finns ett snabbt sätt att utesluta ett visst ord från avstavningen (och rättstavningskontrollen):  
Markera ordet, välj Format - Tecken, klicka på fliken Teckensnitt och välj språket Inget.  
Om du vill utesluta ett ord från den automatiska avstavningen för alltid, så att det aldrig delas, matar du in det med ett likhetstecken efteråt i en aktiverad användarordlista:  
Välj Verktyg - Alternativ - Språkinställningar - Lingvistik  
Välj ut en Användarordlista och klicka på kommandoknappen Redigera.  
Om du inte har någon användarordlista kan du skapa en via kommandoknappen Ny.  
I dialogrutan Redigera användarordlista som öppnas, matar du in ordet t.ex. som "företagsnamn=" (utan citattecknen) och stänger dialogrutorna med Stäng och OK  
Ordet "företagsnamn" avstavas sedan aldrig.  
Du behöver inte söka i texten efter kandidater för manuell avstavning själv.  
Välj kommandot Verktyg - Avstavning.  
Då ser du alla ord, som kan avstavas enligt radbrytningen som gäller, efter varandra i en dialogruta.  
Stället där ordet bäst kan delas vid aktuell radbrytning är markerat.  
Med kommandoknappen Vänsterpil flyttar du markeringen åt vänster om ordet ska delas längre fram.  
När du klickar på Avstava, delas ordet vid markeringen och nästa ord visas som kan avstavas.  
Om ordet är känt i rättstavningskontrollen visas de registrerade avstavningsställena även där.  
Textflöde  
Sätta på / stänga av numreringar  
Så sätter du på och stänger av en numrering  
1.  
Markera styckena som ska numreras.  
2.  
Klicka på ikonen Numrering på / av på textobjektlisten.  
Styckena formateras som numrering.  
Om du klickar på ikonen Numrering på / av i en numrering formateras styckena som normal text igen.  
Det är bäst att ställa in numreringar, precis som punktuppställningar, via ikonerna på Numreringsobjektlisten.  
Om du flyttar en numrering en nivå nedåt börjar numreringen som kommer efter på den här nivån med ett igen.  
De här alternativen finns under Format - Numrering / Punktuppställning - Alternativ.  
Exempel  
1.  
Rad ett  
2. och rad två  
1. och en underordnad nivå till rad 2  
I det här exemplet visas inte numreringen fullständigt.  
Den sista raden med den underordnade nivån till 2. skulle numreras med 2.1. om numreringen var fullständig.  
Sätta på / stänga av punktuppställningar  
Så sätter du på och stänger av en punktuppställning  
1.  
Placera textmarkören i ett stycke som ska markeras med ett punktuppställningstecken eller markera flera stycken.  
2.  
Klicka på ikonen Punktuppställning på / av på textobjektlisten.  
Stycket eller styckena formateras som punktuppställning.  
3.  
Om du klickar på ikonen Punktuppställning på / av i en punktuppställning formateras styckena som normal text igen.  
4.  
I en punktuppställning kan du byta till numreringsobjektlisten med ikonen längst till höger på objektlisten.  
Även på snabbmenyn till objektlisten kan du välja vilken list som ska visas.  
På numreringsobjektlisten finns bl.a. ikoner för att flytta numrerade stycken.  
I dialogrutan Format - Numrering / Punktuppställning kan du göra fler inställningar för den aktuella punktuppställningen där markören finns.  
Om du vill ha ett annat punktuppställningstecken kan du välja det under Format - Numrering / Punktuppställning - Alternativ via kommandoknappen med tre punkter som öppnar dialogrutan Specialtecken.  
Den här kommandoknappen visas bara om du har valt posten "Punkt" i kombinationsfältet Numrering.  
Numrering och numreringsformatmall  
Du kan antingen tilldela numreringarna i dina texter som direkt formatering eller som mall - på samma sätt som andra styckeattribut, t.ex. "Marginaljustering" eller "Radavstånd ".  
Ikonerna på numreringsobjektlisten och alternativen i dialogrutan Format - Numrering / Punktuppställning tilldelar direkta formateringar.  
Även vid automatisk användning av en numrering via AutoFormat / AutoKorrigering-funktionen används direkta formateringar.  
De automatiska numreringarna från AutoKorrigering används inte på mallarna som finns i kategorin "Formatmallar specialområden" i Stylist.  
Du kan tilldela vissa styckeformatmallar en viss Numreringsformatmall eller tilldela styckena numreringsmallen direkt.  
I de här fallen kan du utnyttja fördelarna med mallkonceptet även för numreringar:  
Om du ändrar numreringsformatmallen formateras alla numreringar automatiskt om som du har skapat med den här formatmallen.  
Numreringsformatmallarna beskrivs i %PRODUCTNAME -hjälpen.  
Synonymordlista  
I synonymordlistan kan du slå upp synonymer till ord.  
Markera ordet som du vill hitta synonymer till.  
Välj Verktyg - Synonymordlista eller tryck på Kommando Ctrl +F7.  
En dialogruta öppnas där du kan klicka i de båda undre listrutorna tills du hittar ett lämpligt ord.  
Om du stänger dialogrutan med OK, ersätts det markerade ordet med ordet som står i textfältet Ersätt.  
Synonymordlistan är inte tillgänglig på alla språk för vilka en rättstavningskontroll är installerad.  
Om du letar efter alternativ till ett ord på ett annat språk för vilket en synonymordlista är installerad, t.ex. för ett engelskt ord, markerar du ordet i texten och öppnar synonymordlistan.  
Byt till "Engelska (UK)" eller "Engelska (US) "via kommandoknappen Språk.  
Klicka sedan på Slå upp.  
Om du har givit de engelska orden i din text det engelska språket som attribut (Format - Tecken, fliken Teckensnitt, kombinationsfältet Språk) tar rättstavningskontrollen, synonymordlistan och avstavningen automatiskt hänsyn till det här språket.  
Du kan också tilldela styckeformatmallarna ett språk på motsvarande sätt.  
Synonymordlista  
Räkna ord i text  
Så tar du reda på antalet ord i ett textdokument.  
Under fliken Statistik visas bl.a. antalet använda ord.  
Arkiv - Egenskaper - Statistik  
Textanpassning runt objekt  
Typ av textanpassning kan väljas individuellt för varje objekt.  
Markera objektet och öppna snabbmenyn.  
I snabbmenyn finns de viktigaste alternativen under kommandot Textanpassning.  
Alternativet som gäller i det aktuella fallet är markerat med en punkt i undermenyn.  
Klicka på det textanpassningsalternativ som du vill använda på det markerade objektet.  
Klicka på fliken Textanpassning i dialogrutan.  
De enskilda alternativen beskrivs utförligt i %PRODUCTNAME -hjälpen.  
I den här dialogrutan kan du också ställa in alternativen för formsättningen eller konturanpassningen.  
Om du markerar Kontur kommer texten att följa objektets konturer.  
Om du väljer alternativet Genomflöde anpassas ju inte texten.  
Om du dessutom markerar rutan Bara utanför löper inte texten in i öppna objekt.  
På bilden visas samma objekt med och utan alternativet Bara utanför.  
Du öppnar den via kommandot Textanpassning - Redigera kontur... på snabbmenyn till ett infogat grafikobjekt.  
Den beskrivs utförligt i %PRODUCTNAME -hjälpen.  
Välkommen till %PRODUCTNAME Writer-hjälpen  
Hjälp till %PRODUCTNAME Writer  
Hjälp till hjälpen  
Menyer  
Här finns en beskrivning av alla menyer med undermenyer och dialogrutor som du kan öppna när ett textdokument är aktivt.  
Arkiv  
Du kan t.ex. skapa ett nytt dokument, öppna, stänga och skriva ut dokument, ange dokumentegenskaper med mera.  
När du vill avsluta %PRODUCTNAME klickar du på menykommandot Avsluta.  
Öppna...  
Spara som...  
Versioner...  
Egenskaper...  
Skriv ut...  
Skrivarinställning...  
Kopplad utskrift...  
Redigera  
Här finns även olika funktioner för att redigera förteckningar och integrerade objekt.  
Klistra in innehåll...  
Jämför dokument...  
Sök och ersätt...  
AutoText...  
Byt databas...  
Fältkommando...  
Fotnot...  
Förteckningspost...  
Litteraturförteckningspost  
Hyperlänk  
Länkar...  
Image map  
Visa  
Den här menyn innehåller kommandon som du använder till att styra hur dels %PRODUCTNAME -fönstret ska se ut när ett textdokument är aktivt, dels hur dokumentinnehållet ska se ut på bildskärmen.  
Här kan du bestämma vilka av symbollisterna som ska visas eller i vilken skala du vill att dokumentet ska visas.  
Skala...  
Infoga  
På den här menyn är alla kommandon samlade, som du behöver om du vill infoga nya element i dokumentet, t.ex. områden, fotnoter, anteckningar, extrasidor för kuvert eller etiketter, specialtecken, grafik, objekt från andra tillämpningar o.s.v.  
Manuell brytning...  
Specialtecken...  
Område...  
Hyperlänk  
Fotnot...  
Bildtext...  
Bokmärke...  
Korshänvisning...  
Anteckning...  
Skript  
Kuvert...  
Ram...  
Tabell...  
Horisontell linje...  
Ramteknik  
Fil...  
Format  
Här finns kommandon för textformatering av enskilda tecken, stycken eller hela sidor.  
När andra objekt är markerade, som grafik eller tabeller, ändras menyn så att den innehåller formateringskommandon.  
Om t.ex. grafik är markerad, innehåller formatmenyn bara kommandon som krävs för formatering av grafik, medan kommandona för textformatering inte visas.  
Vidare finns funktionerna för hantering av mallar i den här menyn, t.ex. mallkatalogen och Stylist.  
Tecken...  
Stycke...  
Sida...  
Områden...  
Kolumner...  
Numrering / punktuppställning...  
Följande kommandon visas bara i vissa sammanhang:  
Ram...  
Grafik...  
Objekt...  
Tabell...  
Talformat...  
AutoFormat...  
Linje...  
Yta...  
Text...  
Position och storlek...  
Kontrollfält...  
Formulär...  
Verktyg  
Här startar du rättstavningskontrollen eller synonymordlistan.  
Du styr den automatiska korrigeringen, definierar numrering av kapitel och sidor och mycket annat.  
Du kan också ställa in symbollisternas och menyernas utseende, konfigurera tangentbordet och göra allmänna standardinställningar för programmet.  
Synonymordlista...  
Avstavning...  
AutoKorrigering / AutoFormat...  
Kapitelnumrering...  
Radnumrering...  
Fotnoter...  
Datakällor  
Text <-> Tabell...  
Sortera...  
Makro...  
Anpassa...  
Fönster  
På fönstermenyn kan du öppna nya fönster.  
Här finns även en lista över alla öppna dokument.  
Symbollister  
Här hittar du en beskrivning av hur symbollisterna ser ut när ett textdokumentet är aktivt.  
Textobjektlist  
I textinmatningsläget ser du den här listen med funktioner för formatering av text.  
Här finns de vanligaste funktionerna för direkt teckenformatering, alltså för formatering utan användning av formatmallar.  
Teckenfärg  
Objektlist vid grafik  
Objektlisten innehåller viktiga funktioner för hantering av grafikobjekt.  
Precis som andra symbollister kan du konfigurera den efter dina behov.  
Välj bara menyn Visa - Symbollister - Redigera.  
Spegelvänd vertikalt  
Ikonen motsvarar kryssrutan vertikalt under fliken Grafik.  
Spegelvänd horisontellt  
Ikonen motsvarar kryssrutan horisontalt under fliken Grafik.  
Grafikegenskaper  
Objektlist vid tabeller  
Objektlisten som du får om du placerar markören i en tabell visar de viktigaste funktionerna som du behöver när du arbetar med en tabell, t.ex. infoga och radera rader och kolumner eller ändra linjestil.  
Förbind celler  
Radera rad  
Radera kolumn  
Objektlist vid teckningar  
Om en teckning är markerad innehåller objektlisten de viktigaste funktionerna som du behöver när du ska redigera teckningen, t.ex. linjetjocklek och -färg, placering i för - eller bakgrunden med mera.  
Linjestil  
Linjebredd  
Linjefärg  
Ytstil / -fyllning  
Objektlist vid numreringar  
Med hjälp av objektlisten vid numreringar kan du lätt ändra de numrerade styckenas struktur.  
Du kan sortera om stycken eller definiera olika styckenivåer med ikonerna.  
Statuslisten  
Statuslisten visar information om det aktuella dokumentet och innehåller några kommandoknappar med specialfunktioner.  
Statuslistens visning och funktioner är beroende av vilket objekt du redigerar och vilket fönster som för tillfället är aktivt i arbetsområdet.  
Du kan konfigurera statuslisten precis som andra lister (i dialogrutan under Verktyg - Anpassa...).  
Förhandsgranskning  
Listen med namnet Förhandsgranskning visas om du har aktiverat förhandsgranskningen av det aktuella dokumentet.  
Linjaler  
På linjalerna visas inte bara sidans mått, utan här finns också markeringar för tabbar, indrag, marginaler och kolumner som du kan ändra interaktivt med hjälp av musen.  
Om du dubbelklickar i ett ledigt (grått) område på linjalerna öppnas dialogrutan Stycke där du kan ange direkta styckeformateringar för det aktuella stycket eller alla markerade stycken.  
Formellisten  
Formellisten för textdokument använder du när du vill göra beräkningar.  
Tryck på F2 när du vill aktivera formellisten.  
Objektlist vid ram  
När ramar är markerade innehåller objektlisten de viktigaste funktionerna som du behöver när du ska formatera och justera ramar.  
Textanpassning av  
Den här inställningen kan du också definiera under fliken Textanpassning.  
Textanpassning på  
Vad gäller funktionen motsvarar den här ikonen alternativet Textanpassning sida under fliken Textanpassning.  
Textgenomflöde  
Detta kan du också styra via fliken Textanpassning.  
Bakgrundsfärg  
Ramegenskaper  
Objektlist vid objekt  
När objekt är markerade innehåller objektlisten de viktigaste funktionerna som du behöver till att formatera och justera objekt.  
Textanpassning av  
Den här inställningen kan du också definiera under fliken Textanpassning.  
Textanpassning på  
Vad gäller funktionen motsvarar den här ikonen alternativet Textanpassning sida under fliken Textanpassning.  
Textgenomflöde  
Detta kan du också styra via fliken Textanpassning.  
Objektegenskaper  
Verktygslist  
Med verktygslisten kan du bl.a. infoga objekt av alla slag i dokumentet och snabbt komma åt de mest använda funktionerna.  
Formulär  
Verktygslist / Webb  
Verktygslisten / Webb visas om du har öppnat ett HTML-dokument.  
Du kan infoga objekt av alla slag i dokumentet och snabbt komma åt de mest använda funktionerna.  
Dessutom kan du välja speciella kommandon för HTML-dokument, som t.ex. HTML-källtext.  
Formulär-kontrollfält  
Redigera AutoText  
Objektlist för text i ritobjekt  
Den här objektlisten visas när du placerar textmarkören i ett ritobjekt genom att dubbelklicka så att du kan skriva en text som sitter ihop med objektet.  
Upphöjt  
Nedsänkt  
Markera allt  
Teckenattribut  
Format: stycke  
Här kan du ställa in indrag, avstånd, justering och radavstånd för det markerade stycket.  
Funktioner i %PRODUCTNAME Writer  
Här får du en kort överblick över några viktiga funktioner i %PRODUCTNAME Writer.  
Skriva  
Med %PRODUCTNAME Writer kan du skapa textdokument av alla slag.  
Du kan skapa privatbrev, standardbrev (kopplad utskrift), broschyrer, faxmeddelanden eller professionella handböcker.  
Dokument som du ofta använder kan du spara som mall, t.ex. för ett fakturaformulär.  
Om du vill kan du använda automatisk korrigering och avstavning medan du skriver.  
I %PRODUCTNAME kan du skapa textdokument som kan vara nästan hur långa som helst; med Navigator hittar du ändå snabbt och enkelt dit du vill i dokumentet.  
Med hjälp av AutoPiloterna kan du dessutom enkelt skapa egna skräddarsydda mallar.  
Utforma och strukturera  
Programmet innehåller många möjligheter för att utforma dokument.  
Med Stylist kan du skapa, tilldela och ändra mallar för stycken, tecken, ramar och sidor.  
Med Navigator kan du dessutom snabbt och enkelt göra en disposition av texten och snabbt ändra dispositionen vid behov, t.ex. genom att flytta stycken.  
Du kan då i stor utsträckning själv bestämma hur de ska struktureras och se ut.  
Via hyperlänkar och bokmärken kan du hoppa direkt till ett textställe.  
Desktop Publishing med %PRODUCTNAME Writer  
Du kan sätta texter i flera kolumner och integrera textramar, grafik, tabeller med mera.  
Textramarna kan du länka till varandra kors och tvärs och över sidgränserna som du vill, vilket du har stor nytta av om du vill skapa en tidningslayout.  
Funktioner som radregister, konturflöde runt och genom bilder och valfri färgläggning av tecken, stycken och tabeller gör det ännu lättare att skapa dokument med ett professionellt utseende.  
Göra beräkningar  
I %PRODUCTNAME finns en integrerad räknefunktion för textdokument, med vilken du även kan utföra komplicerade beräkningar eller framställa logiska samband.  
Tabellen som behövs för beräkningar skapar du snabbt och enkelt i textdokumentet.  
Skapa teckningar  
Med hjälp av ett ritverktyg kan du skapa teckningar, grafik, förklaringar och mycket annat direkt i ett textdokument.  
Infoga grafik  
I ett textdokument kan du lägga in grafik i olika format, t.ex. JPG och GIF.  
Det går bra att redigera bilderna direkt i ordbehandlingsdokumentet med programmet för bildredigering.  
Dessutom hittar du ett stort antal clip art-bilder ordnade efter olika teman i Gallery.  
Flexibelt programgränssnitt  
Programgränssnittet är utformat så att alla användare kan konfigurera det individuellt.  
Du kan flytta de olika fönstren (Stylist, Navigator m.fl.) fritt på bildskärmen och delvis kan du förankra dem.  
Dessutom går det att anpassa ikoner och menyer.  
Dra-och-släpp  
Med hjälp av dra-och-släpp (Drag&Drop) kan du arbeta snabbt och intuitivt med textdokument i %PRODUCTNAME.  
Du kan t.ex. dra grafikobjekt direkt från Gallery till det aktuella dokumentet.  
Omfattande hjälpfunktioner  
Programmet har en omfattande hjälpfunktion där det finns en beskrivning av programelementen i %PRODUCTNAME och en mängd anvisningar för både enkla och lite svårare uppgifter.  
